magic
tech scmos
timestamp 1669707107
<< nwell >>
rect -2023 166 -2000 237
rect -1934 165 -1911 236
rect -1847 165 -1824 236
rect -1758 166 -1735 237
rect -1670 166 -1647 237
rect -1580 166 -1557 237
rect -1488 166 -1465 237
rect -1393 166 -1370 237
rect -1304 166 -1281 237
rect -1212 167 -1189 238
rect -1118 166 -1095 237
rect -1030 166 -1007 237
rect -940 166 -917 237
rect -849 166 -826 237
rect -758 166 -735 237
rect -669 166 -646 237
rect -2274 -175 -2214 -4
rect -1986 -97 -1926 74
rect -1769 -39 -1746 32
rect -1696 29 -1673 54
rect -1637 28 -1614 53
rect -1664 -48 -1614 10
rect -1353 -49 -1330 22
rect -1280 19 -1257 44
rect -1221 18 -1198 43
rect -1248 -58 -1198 0
rect -905 -16 -882 55
rect -832 52 -809 77
rect -773 51 -750 76
rect -800 -25 -750 33
rect -2044 -138 -2021 -113
rect -1948 -121 -1926 -97
rect -2332 -216 -2309 -191
rect -2236 -199 -2214 -175
rect -1743 -337 -1683 -166
rect -1492 -297 -1432 -126
rect -1074 -248 -1014 -77
rect -1132 -289 -1109 -264
rect -1036 -272 -1014 -248
rect -2017 -517 -1957 -346
rect -1801 -378 -1778 -353
rect -1705 -361 -1683 -337
rect -1550 -338 -1527 -313
rect -1454 -321 -1432 -297
rect -2075 -558 -2052 -533
rect -1979 -541 -1957 -517
rect -1750 -637 -1690 -466
rect -1601 -536 -1578 -465
rect -1528 -468 -1505 -443
rect -1469 -469 -1446 -444
rect -1291 -484 -1231 -313
rect -1496 -545 -1446 -487
rect -1349 -525 -1326 -500
rect -1253 -508 -1231 -484
rect -1808 -678 -1785 -653
rect -1712 -661 -1690 -637
<< polysilicon >>
rect -2072 220 -2051 222
rect -2072 191 -2070 220
rect -2053 209 -2051 220
rect -2035 219 -2017 221
rect -2009 219 -2005 221
rect -1983 219 -1962 221
rect -2035 209 -2033 219
rect -2063 207 -2060 209
rect -2056 207 -2051 209
rect -2046 207 -2043 209
rect -2039 207 -2033 209
rect -2055 197 -2017 199
rect -2009 197 -2005 199
rect -2055 191 -2053 197
rect -2072 189 -2053 191
rect -1983 190 -1981 219
rect -1964 208 -1962 219
rect -1946 218 -1928 220
rect -1920 218 -1916 220
rect -1896 219 -1875 221
rect -1807 220 -1786 222
rect -1946 208 -1944 218
rect -1974 206 -1971 208
rect -1967 206 -1962 208
rect -1957 206 -1954 208
rect -1950 206 -1944 208
rect -1966 196 -1928 198
rect -1920 196 -1916 198
rect -1966 190 -1964 196
rect -1983 188 -1964 190
rect -1896 190 -1894 219
rect -1877 208 -1875 219
rect -1859 218 -1841 220
rect -1833 218 -1829 220
rect -1859 208 -1857 218
rect -1887 206 -1884 208
rect -1880 206 -1875 208
rect -1870 206 -1867 208
rect -1863 206 -1857 208
rect -1879 196 -1841 198
rect -1833 196 -1829 198
rect -1879 190 -1877 196
rect -1807 191 -1805 220
rect -1788 209 -1786 220
rect -1770 219 -1752 221
rect -1744 219 -1740 221
rect -1719 220 -1698 222
rect -1770 209 -1768 219
rect -1798 207 -1795 209
rect -1791 207 -1786 209
rect -1781 207 -1778 209
rect -1774 207 -1768 209
rect -1790 197 -1752 199
rect -1744 197 -1740 199
rect -1790 191 -1788 197
rect -1896 188 -1877 190
rect -1807 189 -1788 191
rect -1719 191 -1717 220
rect -1700 209 -1698 220
rect -1682 219 -1664 221
rect -1656 219 -1652 221
rect -1629 220 -1608 222
rect -1682 209 -1680 219
rect -1710 207 -1707 209
rect -1703 207 -1698 209
rect -1693 207 -1690 209
rect -1686 207 -1680 209
rect -1702 197 -1664 199
rect -1656 197 -1652 199
rect -1702 191 -1700 197
rect -1719 189 -1700 191
rect -1629 191 -1627 220
rect -1610 209 -1608 220
rect -1592 219 -1574 221
rect -1566 219 -1562 221
rect -1537 220 -1516 222
rect -1592 209 -1590 219
rect -1620 207 -1617 209
rect -1613 207 -1608 209
rect -1603 207 -1600 209
rect -1596 207 -1590 209
rect -1612 197 -1574 199
rect -1566 197 -1562 199
rect -1612 191 -1610 197
rect -1629 189 -1610 191
rect -1537 191 -1535 220
rect -1518 209 -1516 220
rect -1500 219 -1482 221
rect -1474 219 -1470 221
rect -1442 220 -1421 222
rect -1500 209 -1498 219
rect -1528 207 -1525 209
rect -1521 207 -1516 209
rect -1511 207 -1508 209
rect -1504 207 -1498 209
rect -1520 197 -1482 199
rect -1474 197 -1470 199
rect -1520 191 -1518 197
rect -1537 189 -1518 191
rect -1442 191 -1440 220
rect -1423 209 -1421 220
rect -1405 219 -1387 221
rect -1379 219 -1375 221
rect -1353 220 -1332 222
rect -1261 221 -1240 223
rect -1405 209 -1403 219
rect -1433 207 -1430 209
rect -1426 207 -1421 209
rect -1416 207 -1413 209
rect -1409 207 -1403 209
rect -1425 197 -1387 199
rect -1379 197 -1375 199
rect -1425 191 -1423 197
rect -1442 189 -1423 191
rect -1353 191 -1351 220
rect -1334 209 -1332 220
rect -1316 219 -1298 221
rect -1290 219 -1286 221
rect -1316 209 -1314 219
rect -1344 207 -1341 209
rect -1337 207 -1332 209
rect -1327 207 -1324 209
rect -1320 207 -1314 209
rect -1336 197 -1298 199
rect -1290 197 -1286 199
rect -1336 191 -1334 197
rect -1261 192 -1259 221
rect -1242 210 -1240 221
rect -1224 220 -1206 222
rect -1198 220 -1194 222
rect -1167 220 -1146 222
rect -1224 210 -1222 220
rect -1252 208 -1249 210
rect -1245 208 -1240 210
rect -1235 208 -1232 210
rect -1228 208 -1222 210
rect -1244 198 -1206 200
rect -1198 198 -1194 200
rect -1244 192 -1242 198
rect -1353 189 -1334 191
rect -1261 190 -1242 192
rect -1167 191 -1165 220
rect -1148 209 -1146 220
rect -1130 219 -1112 221
rect -1104 219 -1100 221
rect -1079 220 -1058 222
rect -1130 209 -1128 219
rect -1158 207 -1155 209
rect -1151 207 -1146 209
rect -1141 207 -1138 209
rect -1134 207 -1128 209
rect -1150 197 -1112 199
rect -1104 197 -1100 199
rect -1150 191 -1148 197
rect -1167 189 -1148 191
rect -1079 191 -1077 220
rect -1060 209 -1058 220
rect -1042 219 -1024 221
rect -1016 219 -1012 221
rect -989 220 -968 222
rect -1042 209 -1040 219
rect -1070 207 -1067 209
rect -1063 207 -1058 209
rect -1053 207 -1050 209
rect -1046 207 -1040 209
rect -1062 197 -1024 199
rect -1016 197 -1012 199
rect -1062 191 -1060 197
rect -1079 189 -1060 191
rect -989 191 -987 220
rect -970 209 -968 220
rect -952 219 -934 221
rect -926 219 -922 221
rect -898 220 -877 222
rect -952 209 -950 219
rect -980 207 -977 209
rect -973 207 -968 209
rect -963 207 -960 209
rect -956 207 -950 209
rect -972 197 -934 199
rect -926 197 -922 199
rect -972 191 -970 197
rect -989 189 -970 191
rect -898 191 -896 220
rect -879 209 -877 220
rect -861 219 -843 221
rect -835 219 -831 221
rect -807 220 -786 222
rect -861 209 -859 219
rect -889 207 -886 209
rect -882 207 -877 209
rect -872 207 -869 209
rect -865 207 -859 209
rect -881 197 -843 199
rect -835 197 -831 199
rect -881 191 -879 197
rect -898 189 -879 191
rect -807 191 -805 220
rect -788 209 -786 220
rect -770 219 -752 221
rect -744 219 -740 221
rect -718 220 -697 222
rect -770 209 -768 219
rect -798 207 -795 209
rect -791 207 -786 209
rect -781 207 -778 209
rect -774 207 -768 209
rect -790 197 -752 199
rect -744 197 -740 199
rect -790 191 -788 197
rect -807 189 -788 191
rect -718 191 -716 220
rect -699 209 -697 220
rect -681 219 -663 221
rect -655 219 -651 221
rect -681 209 -679 219
rect -709 207 -706 209
rect -702 207 -697 209
rect -692 207 -689 209
rect -685 207 -679 209
rect -701 197 -663 199
rect -655 197 -651 199
rect -701 191 -699 197
rect -718 189 -699 191
rect -2045 178 -2042 180
rect -2038 178 -2017 180
rect -2009 178 -2005 180
rect -1956 177 -1953 179
rect -1949 177 -1928 179
rect -1920 177 -1916 179
rect -1869 177 -1866 179
rect -1862 177 -1841 179
rect -1833 177 -1829 179
rect -1780 178 -1777 180
rect -1773 178 -1752 180
rect -1744 178 -1740 180
rect -1692 178 -1689 180
rect -1685 178 -1664 180
rect -1656 178 -1652 180
rect -1602 178 -1599 180
rect -1595 178 -1574 180
rect -1566 178 -1562 180
rect -1510 178 -1507 180
rect -1503 178 -1482 180
rect -1474 178 -1470 180
rect -1415 178 -1412 180
rect -1408 178 -1387 180
rect -1379 178 -1375 180
rect -1326 178 -1323 180
rect -1319 178 -1298 180
rect -1290 178 -1286 180
rect -1234 179 -1231 181
rect -1227 179 -1206 181
rect -1199 179 -1194 181
rect -1140 178 -1137 180
rect -1133 178 -1112 180
rect -1104 178 -1100 180
rect -1052 178 -1049 180
rect -1045 178 -1024 180
rect -1016 178 -1012 180
rect -962 178 -959 180
rect -955 178 -934 180
rect -926 178 -922 180
rect -871 178 -868 180
rect -864 178 -843 180
rect -835 178 -831 180
rect -780 178 -777 180
rect -773 178 -752 180
rect -744 178 -740 180
rect -691 178 -688 180
rect -684 178 -663 180
rect -655 178 -651 180
rect -2050 71 -1944 73
rect -2050 63 -2048 71
rect -1946 63 -1944 71
rect -851 64 -848 66
rect -844 64 -826 66
rect -818 64 -814 66
rect -2064 61 -2061 63
rect -2057 61 -2048 63
rect -2032 61 -2028 63
rect -2024 61 -1980 63
rect -1972 61 -1969 63
rect -1946 61 -1941 63
rect -1933 61 -1930 63
rect -792 63 -789 65
rect -785 63 -767 65
rect -759 63 -755 65
rect -1715 41 -1712 43
rect -1708 41 -1690 43
rect -1682 41 -1678 43
rect -2065 37 -2061 39
rect -2057 37 -1941 39
rect -1933 37 -1930 39
rect -1656 40 -1653 42
rect -1649 40 -1631 42
rect -1623 40 -1619 42
rect -954 38 -933 40
rect -1299 31 -1296 33
rect -1292 31 -1274 33
rect -1266 31 -1262 33
rect -2032 25 -2028 27
rect -2024 25 -1980 27
rect -1972 25 -1968 27
rect -1240 30 -1237 32
rect -1233 30 -1215 32
rect -1207 30 -1203 32
rect -1818 15 -1797 17
rect -2065 13 -2061 15
rect -2057 13 -1941 15
rect -1933 13 -1930 15
rect -2338 -7 -2232 -5
rect -2338 -15 -2336 -7
rect -2234 -15 -2232 -7
rect -2064 -11 -2061 -9
rect -2057 -11 -1941 -9
rect -1933 -11 -1930 -9
rect -2352 -17 -2349 -15
rect -2345 -17 -2336 -15
rect -2320 -17 -2316 -15
rect -2312 -17 -2268 -15
rect -2260 -17 -2257 -15
rect -2234 -17 -2229 -15
rect -2221 -17 -2218 -15
rect -1818 -14 -1816 15
rect -1799 4 -1797 15
rect -1781 14 -1763 16
rect -1755 14 -1751 16
rect -1781 4 -1779 14
rect -1701 13 -1675 15
rect -1809 2 -1806 4
rect -1802 2 -1797 4
rect -1792 2 -1789 4
rect -1785 2 -1779 4
rect -1701 -2 -1699 13
rect -1677 -1 -1675 13
rect -1402 5 -1381 7
rect -954 9 -952 38
rect -935 27 -933 38
rect -917 37 -899 39
rect -891 37 -887 39
rect -917 27 -915 37
rect -837 36 -811 38
rect -945 25 -942 27
rect -938 25 -933 27
rect -928 25 -925 27
rect -921 25 -915 27
rect -837 21 -835 36
rect -813 22 -811 36
rect -848 19 -845 21
rect -841 19 -835 21
rect -827 20 -823 22
rect -819 20 -816 22
rect -813 20 -794 22
rect -786 20 -781 22
rect -772 20 -768 22
rect -760 20 -757 22
rect -937 15 -899 17
rect -891 15 -887 17
rect -937 9 -935 15
rect -954 7 -935 9
rect -1712 -4 -1709 -2
rect -1705 -4 -1699 -2
rect -1691 -3 -1687 -1
rect -1683 -3 -1680 -1
rect -1677 -3 -1658 -1
rect -1650 -3 -1645 -1
rect -1636 -3 -1632 -1
rect -1624 -3 -1621 -1
rect -1801 -8 -1763 -6
rect -1755 -8 -1751 -6
rect -1801 -14 -1799 -8
rect -1818 -16 -1799 -14
rect -1691 -18 -1689 -3
rect -1722 -20 -1689 -18
rect -1791 -27 -1788 -25
rect -1784 -27 -1763 -25
rect -1755 -27 -1751 -25
rect -2064 -35 -2061 -33
rect -2057 -35 -2044 -33
rect -2032 -35 -2028 -33
rect -2024 -35 -1980 -33
rect -1972 -35 -1967 -33
rect -1951 -35 -1941 -33
rect -1933 -35 -1930 -33
rect -2353 -41 -2349 -39
rect -2345 -41 -2229 -39
rect -2221 -41 -2218 -39
rect -2046 -44 -2044 -35
rect -1951 -44 -1949 -35
rect -2046 -46 -1949 -44
rect -2320 -53 -2316 -51
rect -2312 -53 -2268 -51
rect -2260 -53 -2256 -51
rect -2064 -59 -2061 -57
rect -2057 -59 -1941 -57
rect -1933 -59 -1930 -57
rect -2353 -65 -2349 -63
rect -2345 -65 -2229 -63
rect -2221 -65 -2218 -63
rect -1722 -66 -1720 -20
rect -1636 -26 -1634 -3
rect -1402 -24 -1400 5
rect -1383 -6 -1381 5
rect -1365 4 -1347 6
rect -1339 4 -1335 6
rect -827 5 -825 20
rect -1365 -6 -1363 4
rect -1285 3 -1259 5
rect -858 3 -825 5
rect -1393 -8 -1390 -6
rect -1386 -8 -1381 -6
rect -1376 -8 -1373 -6
rect -1369 -8 -1363 -6
rect -1285 -12 -1283 3
rect -1261 -11 -1259 3
rect -927 -4 -924 -2
rect -920 -4 -899 -2
rect -891 -4 -887 -2
rect -1296 -14 -1293 -12
rect -1289 -14 -1283 -12
rect -1275 -13 -1271 -11
rect -1267 -13 -1264 -11
rect -1261 -13 -1242 -11
rect -1234 -13 -1229 -11
rect -1220 -13 -1216 -11
rect -1208 -13 -1205 -11
rect -1385 -18 -1347 -16
rect -1339 -18 -1335 -16
rect -1385 -24 -1383 -18
rect -1402 -26 -1383 -24
rect -1672 -28 -1634 -26
rect -1275 -28 -1273 -13
rect -1712 -31 -1709 -29
rect -1705 -31 -1699 -29
rect -1691 -30 -1687 -28
rect -1683 -30 -1670 -28
rect -1306 -30 -1273 -28
rect -1701 -47 -1699 -31
rect -1670 -37 -1658 -35
rect -1650 -37 -1646 -35
rect -1636 -37 -1632 -35
rect -1624 -37 -1621 -35
rect -1375 -37 -1372 -35
rect -1368 -37 -1347 -35
rect -1339 -37 -1335 -35
rect -1670 -47 -1668 -37
rect -1701 -49 -1668 -47
rect -1636 -66 -1634 -37
rect -1722 -68 -1634 -66
rect -2055 -73 -1942 -71
rect -2055 -81 -2053 -73
rect -1944 -81 -1942 -73
rect -1306 -76 -1304 -30
rect -1220 -36 -1218 -13
rect -1256 -38 -1218 -36
rect -1296 -41 -1293 -39
rect -1289 -41 -1283 -39
rect -1275 -40 -1271 -38
rect -1267 -40 -1254 -38
rect -1285 -57 -1283 -41
rect -858 -43 -856 3
rect -772 -3 -770 20
rect -808 -5 -770 -3
rect -848 -8 -845 -6
rect -841 -8 -835 -6
rect -827 -7 -823 -5
rect -819 -7 -806 -5
rect -837 -24 -835 -8
rect -806 -14 -794 -12
rect -786 -14 -782 -12
rect -772 -14 -768 -12
rect -760 -14 -757 -12
rect -806 -24 -804 -14
rect -837 -26 -804 -24
rect -772 -43 -770 -14
rect -858 -45 -770 -43
rect -1254 -47 -1242 -45
rect -1234 -47 -1230 -45
rect -1220 -47 -1216 -45
rect -1208 -47 -1205 -45
rect -1254 -57 -1252 -47
rect -1285 -59 -1252 -57
rect -1220 -76 -1218 -47
rect -1306 -78 -1218 -76
rect -1138 -80 -1032 -78
rect -2064 -83 -2061 -81
rect -2057 -83 -2053 -81
rect -2047 -83 -2044 -81
rect -2040 -83 -2037 -81
rect -2030 -83 -2028 -81
rect -2024 -83 -1980 -81
rect -1972 -83 -1970 -81
rect -1964 -83 -1961 -81
rect -1953 -83 -1949 -81
rect -1944 -83 -1941 -81
rect -1933 -83 -1930 -81
rect -2352 -89 -2349 -87
rect -2345 -89 -2229 -87
rect -2221 -89 -2218 -87
rect -2039 -93 -2037 -83
rect -1964 -93 -1962 -83
rect -1138 -88 -1136 -80
rect -1034 -88 -1032 -80
rect -1152 -90 -1149 -88
rect -1145 -90 -1136 -88
rect -1120 -90 -1116 -88
rect -1112 -90 -1068 -88
rect -1060 -90 -1057 -88
rect -1034 -90 -1029 -88
rect -1021 -90 -1018 -88
rect -2039 -95 -1962 -93
rect -1972 -111 -1968 -109
rect -1964 -111 -1941 -109
rect -1933 -111 -1930 -109
rect -2352 -113 -2349 -111
rect -2345 -113 -2332 -111
rect -2320 -113 -2316 -111
rect -2312 -113 -2268 -111
rect -2260 -113 -2255 -111
rect -2239 -113 -2229 -111
rect -2221 -113 -2218 -111
rect -2334 -122 -2332 -113
rect -2239 -122 -2237 -113
rect -1153 -114 -1149 -112
rect -1145 -114 -1029 -112
rect -1021 -114 -1018 -112
rect -2334 -124 -2237 -122
rect -2065 -126 -2061 -124
rect -2057 -126 -2036 -124
rect -2028 -126 -2024 -124
rect -1120 -126 -1116 -124
rect -1112 -126 -1068 -124
rect -1060 -126 -1056 -124
rect -1556 -129 -1450 -127
rect -2352 -137 -2349 -135
rect -2345 -137 -2229 -135
rect -2221 -137 -2218 -135
rect -1556 -137 -1554 -129
rect -1452 -137 -1450 -129
rect -1570 -139 -1567 -137
rect -1563 -139 -1554 -137
rect -1538 -139 -1534 -137
rect -1530 -139 -1486 -137
rect -1478 -139 -1475 -137
rect -1452 -139 -1447 -137
rect -1439 -139 -1436 -137
rect -1153 -138 -1149 -136
rect -1145 -138 -1029 -136
rect -1021 -138 -1018 -136
rect -2343 -151 -2230 -149
rect -2343 -159 -2341 -151
rect -2232 -159 -2230 -151
rect -2352 -161 -2349 -159
rect -2345 -161 -2341 -159
rect -2335 -161 -2332 -159
rect -2328 -161 -2325 -159
rect -2318 -161 -2316 -159
rect -2312 -161 -2268 -159
rect -2260 -161 -2258 -159
rect -2252 -161 -2249 -159
rect -2241 -161 -2237 -159
rect -2232 -161 -2229 -159
rect -2221 -161 -2218 -159
rect -2327 -171 -2325 -161
rect -2252 -171 -2250 -161
rect -1571 -163 -1567 -161
rect -1563 -163 -1447 -161
rect -1439 -163 -1436 -161
rect -1152 -162 -1149 -160
rect -1145 -162 -1029 -160
rect -1021 -162 -1018 -160
rect -1807 -169 -1701 -167
rect -2327 -173 -2250 -171
rect -1807 -177 -1805 -169
rect -1703 -177 -1701 -169
rect -1538 -175 -1534 -173
rect -1530 -175 -1486 -173
rect -1478 -175 -1474 -173
rect -1821 -179 -1818 -177
rect -1814 -179 -1805 -177
rect -1789 -179 -1785 -177
rect -1781 -179 -1737 -177
rect -1729 -179 -1726 -177
rect -1703 -179 -1698 -177
rect -1690 -179 -1687 -177
rect -1571 -187 -1567 -185
rect -1563 -187 -1447 -185
rect -1439 -187 -1436 -185
rect -1152 -186 -1149 -184
rect -1145 -186 -1132 -184
rect -1120 -186 -1116 -184
rect -1112 -186 -1068 -184
rect -1060 -186 -1055 -184
rect -1039 -186 -1029 -184
rect -1021 -186 -1018 -184
rect -2260 -189 -2256 -187
rect -2252 -189 -2229 -187
rect -2221 -189 -2218 -187
rect -1134 -195 -1132 -186
rect -1039 -195 -1037 -186
rect -1134 -197 -1037 -195
rect -2353 -204 -2349 -202
rect -2345 -204 -2324 -202
rect -2316 -204 -2312 -202
rect -1822 -203 -1818 -201
rect -1814 -203 -1698 -201
rect -1690 -203 -1687 -201
rect -1570 -211 -1567 -209
rect -1563 -211 -1447 -209
rect -1439 -211 -1436 -209
rect -1152 -210 -1149 -208
rect -1145 -210 -1029 -208
rect -1021 -210 -1018 -208
rect -1789 -215 -1785 -213
rect -1781 -215 -1737 -213
rect -1729 -215 -1725 -213
rect -1143 -224 -1030 -222
rect -1822 -227 -1818 -225
rect -1814 -227 -1698 -225
rect -1690 -227 -1687 -225
rect -1143 -232 -1141 -224
rect -1032 -232 -1030 -224
rect -1570 -235 -1567 -233
rect -1563 -235 -1550 -233
rect -1538 -235 -1534 -233
rect -1530 -235 -1486 -233
rect -1478 -235 -1473 -233
rect -1457 -235 -1447 -233
rect -1439 -235 -1436 -233
rect -1152 -234 -1149 -232
rect -1145 -234 -1141 -232
rect -1135 -234 -1132 -232
rect -1128 -234 -1125 -232
rect -1118 -234 -1116 -232
rect -1112 -234 -1068 -232
rect -1060 -234 -1058 -232
rect -1052 -234 -1049 -232
rect -1041 -234 -1037 -232
rect -1032 -234 -1029 -232
rect -1021 -234 -1018 -232
rect -1552 -244 -1550 -235
rect -1457 -244 -1455 -235
rect -1552 -246 -1455 -244
rect -1127 -244 -1125 -234
rect -1052 -244 -1050 -234
rect -1127 -246 -1050 -244
rect -1821 -251 -1818 -249
rect -1814 -251 -1698 -249
rect -1690 -251 -1687 -249
rect -1570 -259 -1567 -257
rect -1563 -259 -1447 -257
rect -1439 -259 -1436 -257
rect -1060 -262 -1056 -260
rect -1052 -262 -1029 -260
rect -1021 -262 -1018 -260
rect -1561 -273 -1448 -271
rect -1821 -275 -1818 -273
rect -1814 -275 -1801 -273
rect -1789 -275 -1785 -273
rect -1781 -275 -1737 -273
rect -1729 -275 -1724 -273
rect -1708 -275 -1698 -273
rect -1690 -275 -1687 -273
rect -1803 -284 -1801 -275
rect -1708 -284 -1706 -275
rect -1561 -281 -1559 -273
rect -1450 -281 -1448 -273
rect -1153 -277 -1149 -275
rect -1145 -277 -1124 -275
rect -1116 -277 -1112 -275
rect -1570 -283 -1567 -281
rect -1563 -283 -1559 -281
rect -1553 -283 -1550 -281
rect -1546 -283 -1543 -281
rect -1536 -283 -1534 -281
rect -1530 -283 -1486 -281
rect -1478 -283 -1476 -281
rect -1470 -283 -1467 -281
rect -1459 -283 -1455 -281
rect -1450 -283 -1447 -281
rect -1439 -283 -1436 -281
rect -1803 -286 -1706 -284
rect -1545 -293 -1543 -283
rect -1470 -293 -1468 -283
rect -1545 -295 -1468 -293
rect -1821 -299 -1818 -297
rect -1814 -299 -1698 -297
rect -1690 -299 -1687 -297
rect -1478 -311 -1474 -309
rect -1470 -311 -1447 -309
rect -1439 -311 -1436 -309
rect -1812 -313 -1699 -311
rect -1812 -321 -1810 -313
rect -1701 -321 -1699 -313
rect -1355 -316 -1249 -314
rect -1821 -323 -1818 -321
rect -1814 -323 -1810 -321
rect -1804 -323 -1801 -321
rect -1797 -323 -1794 -321
rect -1787 -323 -1785 -321
rect -1781 -323 -1737 -321
rect -1729 -323 -1727 -321
rect -1721 -323 -1718 -321
rect -1710 -323 -1706 -321
rect -1701 -323 -1698 -321
rect -1690 -323 -1687 -321
rect -1796 -333 -1794 -323
rect -1721 -333 -1719 -323
rect -1355 -324 -1353 -316
rect -1251 -324 -1249 -316
rect -1571 -326 -1567 -324
rect -1563 -326 -1542 -324
rect -1534 -326 -1530 -324
rect -1369 -326 -1366 -324
rect -1362 -326 -1353 -324
rect -1337 -326 -1333 -324
rect -1329 -326 -1285 -324
rect -1277 -326 -1274 -324
rect -1251 -326 -1246 -324
rect -1238 -326 -1235 -324
rect -1796 -335 -1719 -333
rect -2081 -349 -1975 -347
rect -2081 -357 -2079 -349
rect -1977 -357 -1975 -349
rect -1729 -351 -1725 -349
rect -1721 -351 -1698 -349
rect -1690 -351 -1687 -349
rect -1370 -350 -1366 -348
rect -1362 -350 -1246 -348
rect -1238 -350 -1235 -348
rect -2095 -359 -2092 -357
rect -2088 -359 -2079 -357
rect -2063 -359 -2059 -357
rect -2055 -359 -2011 -357
rect -2003 -359 -2000 -357
rect -1977 -359 -1972 -357
rect -1964 -359 -1961 -357
rect -1337 -362 -1333 -360
rect -1329 -362 -1285 -360
rect -1277 -362 -1273 -360
rect -1822 -366 -1818 -364
rect -1814 -366 -1793 -364
rect -1785 -366 -1781 -364
rect -1370 -374 -1366 -372
rect -1362 -374 -1246 -372
rect -1238 -374 -1235 -372
rect -2096 -383 -2092 -381
rect -2088 -383 -1972 -381
rect -1964 -383 -1961 -381
rect -2063 -395 -2059 -393
rect -2055 -395 -2011 -393
rect -2003 -395 -1999 -393
rect -1369 -398 -1366 -396
rect -1362 -398 -1246 -396
rect -1238 -398 -1235 -396
rect -2096 -407 -2092 -405
rect -2088 -407 -1972 -405
rect -1964 -407 -1961 -405
rect -1369 -422 -1366 -420
rect -1362 -422 -1349 -420
rect -1337 -422 -1333 -420
rect -1329 -422 -1285 -420
rect -1277 -422 -1272 -420
rect -1256 -422 -1246 -420
rect -1238 -422 -1235 -420
rect -2095 -431 -2092 -429
rect -2088 -431 -1972 -429
rect -1964 -431 -1961 -429
rect -1351 -431 -1349 -422
rect -1256 -431 -1254 -422
rect -1351 -433 -1254 -431
rect -1369 -446 -1366 -444
rect -1362 -446 -1246 -444
rect -1238 -446 -1235 -444
rect -2095 -455 -2092 -453
rect -2088 -455 -2075 -453
rect -2063 -455 -2059 -453
rect -2055 -455 -2011 -453
rect -2003 -455 -1998 -453
rect -1982 -455 -1972 -453
rect -1964 -455 -1961 -453
rect -2077 -464 -2075 -455
rect -1982 -464 -1980 -455
rect -1547 -456 -1544 -454
rect -1540 -456 -1522 -454
rect -1514 -456 -1510 -454
rect -1488 -457 -1485 -455
rect -1481 -457 -1463 -455
rect -1455 -457 -1451 -455
rect -1360 -460 -1247 -458
rect -2077 -466 -1980 -464
rect -1814 -469 -1708 -467
rect -1360 -468 -1358 -460
rect -1249 -468 -1247 -460
rect -1814 -477 -1812 -469
rect -1710 -477 -1708 -469
rect -1369 -470 -1366 -468
rect -1362 -470 -1358 -468
rect -1352 -470 -1349 -468
rect -1345 -470 -1342 -468
rect -1335 -470 -1333 -468
rect -1329 -470 -1285 -468
rect -1277 -470 -1275 -468
rect -1269 -470 -1266 -468
rect -1258 -470 -1254 -468
rect -1249 -470 -1246 -468
rect -1238 -470 -1235 -468
rect -2095 -479 -2092 -477
rect -2088 -479 -1972 -477
rect -1964 -479 -1961 -477
rect -1828 -479 -1825 -477
rect -1821 -479 -1812 -477
rect -1796 -479 -1792 -477
rect -1788 -479 -1744 -477
rect -1736 -479 -1733 -477
rect -1710 -479 -1705 -477
rect -1697 -479 -1694 -477
rect -1650 -482 -1629 -480
rect -1344 -480 -1342 -470
rect -1269 -480 -1267 -470
rect -2086 -493 -1973 -491
rect -2086 -501 -2084 -493
rect -1975 -501 -1973 -493
rect -2095 -503 -2092 -501
rect -2088 -503 -2084 -501
rect -2078 -503 -2075 -501
rect -2071 -503 -2068 -501
rect -2061 -503 -2059 -501
rect -2055 -503 -2011 -501
rect -2003 -503 -2001 -501
rect -1995 -503 -1992 -501
rect -1984 -503 -1980 -501
rect -1975 -503 -1972 -501
rect -1964 -503 -1961 -501
rect -1829 -503 -1825 -501
rect -1821 -503 -1705 -501
rect -1697 -503 -1694 -501
rect -2070 -513 -2068 -503
rect -1995 -513 -1993 -503
rect -2070 -515 -1993 -513
rect -1650 -511 -1648 -482
rect -1631 -493 -1629 -482
rect -1613 -483 -1595 -481
rect -1587 -483 -1583 -481
rect -1344 -482 -1267 -480
rect -1613 -493 -1611 -483
rect -1533 -484 -1507 -482
rect -1641 -495 -1638 -493
rect -1634 -495 -1629 -493
rect -1624 -495 -1621 -493
rect -1617 -495 -1611 -493
rect -1533 -499 -1531 -484
rect -1509 -498 -1507 -484
rect -1277 -498 -1273 -496
rect -1269 -498 -1246 -496
rect -1238 -498 -1235 -496
rect -1544 -501 -1541 -499
rect -1537 -501 -1531 -499
rect -1523 -500 -1519 -498
rect -1515 -500 -1512 -498
rect -1509 -500 -1490 -498
rect -1482 -500 -1477 -498
rect -1468 -500 -1464 -498
rect -1456 -500 -1453 -498
rect -1633 -505 -1595 -503
rect -1587 -505 -1583 -503
rect -1633 -511 -1631 -505
rect -1650 -513 -1631 -511
rect -1796 -515 -1792 -513
rect -1788 -515 -1744 -513
rect -1736 -515 -1732 -513
rect -1523 -515 -1521 -500
rect -1554 -517 -1521 -515
rect -1623 -524 -1620 -522
rect -1616 -524 -1595 -522
rect -1587 -524 -1583 -522
rect -1829 -527 -1825 -525
rect -1821 -527 -1705 -525
rect -1697 -527 -1694 -525
rect -2003 -531 -1999 -529
rect -1995 -531 -1972 -529
rect -1964 -531 -1961 -529
rect -2096 -546 -2092 -544
rect -2088 -546 -2067 -544
rect -2059 -546 -2055 -544
rect -1828 -551 -1825 -549
rect -1821 -551 -1705 -549
rect -1697 -551 -1694 -549
rect -1554 -563 -1552 -517
rect -1468 -523 -1466 -500
rect -1370 -513 -1366 -511
rect -1362 -513 -1341 -511
rect -1333 -513 -1329 -511
rect -1504 -525 -1466 -523
rect -1544 -528 -1541 -526
rect -1537 -528 -1531 -526
rect -1523 -527 -1519 -525
rect -1515 -527 -1502 -525
rect -1533 -544 -1531 -528
rect -1502 -534 -1490 -532
rect -1482 -534 -1478 -532
rect -1468 -534 -1464 -532
rect -1456 -534 -1453 -532
rect -1502 -544 -1500 -534
rect -1533 -546 -1500 -544
rect -1468 -563 -1466 -534
rect -1554 -565 -1466 -563
rect -1828 -575 -1825 -573
rect -1821 -575 -1808 -573
rect -1796 -575 -1792 -573
rect -1788 -575 -1744 -573
rect -1736 -575 -1731 -573
rect -1715 -575 -1705 -573
rect -1697 -575 -1694 -573
rect -1810 -584 -1808 -575
rect -1715 -584 -1713 -575
rect -1810 -586 -1713 -584
rect -1828 -599 -1825 -597
rect -1821 -599 -1705 -597
rect -1697 -599 -1694 -597
rect -1819 -613 -1706 -611
rect -1819 -621 -1817 -613
rect -1708 -621 -1706 -613
rect -1828 -623 -1825 -621
rect -1821 -623 -1817 -621
rect -1811 -623 -1808 -621
rect -1804 -623 -1801 -621
rect -1794 -623 -1792 -621
rect -1788 -623 -1744 -621
rect -1736 -623 -1734 -621
rect -1728 -623 -1725 -621
rect -1717 -623 -1713 -621
rect -1708 -623 -1705 -621
rect -1697 -623 -1694 -621
rect -1803 -633 -1801 -623
rect -1728 -633 -1726 -623
rect -1803 -635 -1726 -633
rect -1736 -651 -1732 -649
rect -1728 -651 -1705 -649
rect -1697 -651 -1694 -649
rect -1829 -666 -1825 -664
rect -1821 -666 -1800 -664
rect -1792 -666 -1788 -664
<< ndiffusion >>
rect -2060 209 -2056 210
rect -2043 209 -2039 210
rect -2060 206 -2056 207
rect -2043 206 -2039 207
rect -1971 208 -1967 209
rect -1954 208 -1950 209
rect -1971 205 -1967 206
rect -1954 205 -1950 206
rect -1884 208 -1880 209
rect -1867 208 -1863 209
rect -1884 205 -1880 206
rect -1867 205 -1863 206
rect -1795 209 -1791 210
rect -1778 209 -1774 210
rect -1795 206 -1791 207
rect -1778 206 -1774 207
rect -1707 209 -1703 210
rect -1690 209 -1686 210
rect -1707 206 -1703 207
rect -1690 206 -1686 207
rect -1617 209 -1613 210
rect -1600 209 -1596 210
rect -1617 206 -1613 207
rect -1600 206 -1596 207
rect -1525 209 -1521 210
rect -1508 209 -1504 210
rect -1525 206 -1521 207
rect -1508 206 -1504 207
rect -1430 209 -1426 210
rect -1413 209 -1409 210
rect -1430 206 -1426 207
rect -1413 206 -1409 207
rect -1341 209 -1337 210
rect -1324 209 -1320 210
rect -1341 206 -1337 207
rect -1324 206 -1320 207
rect -1249 210 -1245 211
rect -1232 210 -1228 211
rect -1249 207 -1245 208
rect -1232 207 -1228 208
rect -1155 209 -1151 210
rect -1138 209 -1134 210
rect -1155 206 -1151 207
rect -1138 206 -1134 207
rect -1067 209 -1063 210
rect -1050 209 -1046 210
rect -1067 206 -1063 207
rect -1050 206 -1046 207
rect -977 209 -973 210
rect -960 209 -956 210
rect -977 206 -973 207
rect -960 206 -956 207
rect -886 209 -882 210
rect -869 209 -865 210
rect -886 206 -882 207
rect -869 206 -865 207
rect -795 209 -791 210
rect -778 209 -774 210
rect -795 206 -791 207
rect -778 206 -774 207
rect -706 209 -702 210
rect -689 209 -685 210
rect -706 206 -702 207
rect -689 206 -685 207
rect -2042 180 -2038 181
rect -1953 179 -1949 180
rect -1866 179 -1862 180
rect -1777 180 -1773 181
rect -1689 180 -1685 181
rect -1599 180 -1595 181
rect -1507 180 -1503 181
rect -1412 180 -1408 181
rect -1323 180 -1319 181
rect -1231 181 -1227 182
rect -2042 177 -2038 178
rect -1137 180 -1133 181
rect -1049 180 -1045 181
rect -959 180 -955 181
rect -868 180 -864 181
rect -777 180 -773 181
rect -688 180 -684 181
rect -1231 178 -1227 179
rect -1777 177 -1773 178
rect -1953 176 -1949 177
rect -1866 176 -1862 177
rect -1689 177 -1685 178
rect -1599 177 -1595 178
rect -1507 177 -1503 178
rect -1412 177 -1408 178
rect -1323 177 -1319 178
rect -1137 177 -1133 178
rect -1049 177 -1045 178
rect -959 177 -955 178
rect -868 177 -864 178
rect -777 177 -773 178
rect -688 177 -684 178
rect -2061 63 -2057 64
rect -2028 63 -2024 64
rect -848 66 -844 67
rect -789 65 -785 70
rect -848 63 -844 64
rect -2061 60 -2057 61
rect -2028 60 -2024 61
rect -789 62 -785 63
rect -2061 39 -2057 40
rect -1712 43 -1708 44
rect -1653 42 -1649 47
rect -1712 40 -1708 41
rect -2061 36 -2057 37
rect -1653 39 -1649 40
rect -1296 33 -1292 34
rect -2028 27 -2024 28
rect -1237 32 -1233 37
rect -1296 30 -1292 31
rect -1237 29 -1233 30
rect -2028 24 -2024 25
rect -2061 15 -2057 16
rect -2061 12 -2057 13
rect -2349 -15 -2345 -14
rect -2316 -15 -2312 -14
rect -2061 -9 -2057 -8
rect -2061 -12 -2057 -11
rect -1806 4 -1802 5
rect -1789 4 -1785 5
rect -1806 1 -1802 2
rect -1789 1 -1785 2
rect -1709 -2 -1705 -1
rect -1687 -1 -1683 0
rect -942 27 -938 28
rect -925 27 -921 28
rect -942 24 -938 25
rect -925 24 -921 25
rect -845 21 -841 22
rect -823 22 -819 23
rect -845 18 -841 19
rect -1709 -5 -1705 -4
rect -2349 -18 -2345 -17
rect -2316 -18 -2312 -17
rect -1687 -4 -1683 -3
rect -1788 -25 -1784 -24
rect -1788 -28 -1784 -27
rect -2061 -33 -2057 -32
rect -2028 -33 -2024 -32
rect -2349 -39 -2345 -38
rect -2061 -36 -2057 -35
rect -2349 -42 -2345 -41
rect -2028 -36 -2024 -35
rect -2316 -51 -2312 -50
rect -2316 -54 -2312 -53
rect -2061 -57 -2057 -56
rect -2349 -63 -2345 -62
rect -2061 -60 -2057 -59
rect -2349 -66 -2345 -65
rect -1390 -6 -1386 -5
rect -823 19 -819 20
rect -1373 -6 -1369 -5
rect -1390 -9 -1386 -8
rect -1373 -9 -1369 -8
rect -1293 -12 -1289 -11
rect -1271 -11 -1267 -10
rect -924 -2 -920 -1
rect -924 -5 -920 -4
rect -1293 -15 -1289 -14
rect -1687 -28 -1683 -27
rect -1271 -14 -1267 -13
rect -1709 -29 -1705 -28
rect -1709 -32 -1705 -31
rect -1687 -31 -1683 -30
rect -1372 -35 -1368 -34
rect -1372 -38 -1368 -37
rect -2061 -81 -2057 -80
rect -2044 -81 -2040 -80
rect -2028 -81 -2024 -80
rect -1271 -38 -1267 -37
rect -1293 -39 -1289 -38
rect -1293 -42 -1289 -41
rect -1271 -41 -1267 -40
rect -823 -5 -819 -4
rect -845 -6 -841 -5
rect -845 -9 -841 -8
rect -823 -8 -819 -7
rect -2349 -87 -2345 -86
rect -2061 -84 -2057 -83
rect -2044 -84 -2040 -83
rect -2349 -90 -2345 -89
rect -2028 -84 -2024 -83
rect -1149 -88 -1145 -87
rect -1116 -88 -1112 -87
rect -1149 -91 -1145 -90
rect -1116 -91 -1112 -90
rect -2349 -111 -2345 -110
rect -2316 -111 -2312 -110
rect -1968 -109 -1964 -108
rect -1968 -112 -1964 -111
rect -2349 -114 -2345 -113
rect -2316 -114 -2312 -113
rect -1149 -112 -1145 -111
rect -1149 -115 -1145 -114
rect -2061 -124 -2057 -123
rect -2061 -127 -2057 -126
rect -2349 -135 -2345 -134
rect -1116 -124 -1112 -123
rect -1116 -127 -1112 -126
rect -1567 -137 -1563 -136
rect -1534 -137 -1530 -136
rect -1149 -136 -1145 -135
rect -2349 -138 -2345 -137
rect -1149 -139 -1145 -138
rect -1567 -140 -1563 -139
rect -1534 -140 -1530 -139
rect -2349 -159 -2345 -158
rect -2332 -159 -2328 -158
rect -2316 -159 -2312 -158
rect -1567 -161 -1563 -160
rect -1149 -160 -1145 -159
rect -2349 -162 -2345 -161
rect -2332 -162 -2328 -161
rect -2316 -162 -2312 -161
rect -1149 -163 -1145 -162
rect -1567 -164 -1563 -163
rect -1818 -177 -1814 -176
rect -1785 -177 -1781 -176
rect -1534 -173 -1530 -172
rect -1534 -176 -1530 -175
rect -1818 -180 -1814 -179
rect -2256 -187 -2252 -186
rect -1785 -180 -1781 -179
rect -1567 -185 -1563 -184
rect -1149 -184 -1145 -183
rect -1116 -184 -1112 -183
rect -1149 -187 -1145 -186
rect -1567 -188 -1563 -187
rect -2256 -190 -2252 -189
rect -1116 -187 -1112 -186
rect -2349 -202 -2345 -201
rect -1818 -201 -1814 -200
rect -1818 -204 -1814 -203
rect -2349 -205 -2345 -204
rect -1785 -213 -1781 -212
rect -1567 -209 -1563 -208
rect -1149 -208 -1145 -207
rect -1149 -211 -1145 -210
rect -1567 -212 -1563 -211
rect -1785 -216 -1781 -215
rect -1818 -225 -1814 -224
rect -1818 -228 -1814 -227
rect -1567 -233 -1563 -232
rect -1534 -233 -1530 -232
rect -1149 -232 -1145 -231
rect -1132 -232 -1128 -231
rect -1116 -232 -1112 -231
rect -1149 -235 -1145 -234
rect -1567 -236 -1563 -235
rect -1534 -236 -1530 -235
rect -1132 -235 -1128 -234
rect -1818 -249 -1814 -248
rect -1116 -235 -1112 -234
rect -1818 -252 -1814 -251
rect -1567 -257 -1563 -256
rect -1567 -260 -1563 -259
rect -1056 -260 -1052 -259
rect -1056 -263 -1052 -262
rect -1818 -273 -1814 -272
rect -1785 -273 -1781 -272
rect -1818 -276 -1814 -275
rect -1785 -276 -1781 -275
rect -1567 -281 -1563 -280
rect -1550 -281 -1546 -280
rect -1534 -281 -1530 -280
rect -1149 -275 -1145 -274
rect -1149 -278 -1145 -277
rect -1567 -284 -1563 -283
rect -1550 -284 -1546 -283
rect -1818 -297 -1814 -296
rect -1534 -284 -1530 -283
rect -1818 -300 -1814 -299
rect -1474 -309 -1470 -308
rect -1818 -321 -1814 -320
rect -1801 -321 -1797 -320
rect -1785 -321 -1781 -320
rect -1474 -312 -1470 -311
rect -1818 -324 -1814 -323
rect -1801 -324 -1797 -323
rect -1785 -324 -1781 -323
rect -1567 -324 -1563 -323
rect -1366 -324 -1362 -323
rect -1333 -324 -1329 -323
rect -1567 -327 -1563 -326
rect -1366 -327 -1362 -326
rect -1333 -327 -1329 -326
rect -1725 -349 -1721 -348
rect -1366 -348 -1362 -347
rect -2092 -357 -2088 -356
rect -2059 -357 -2055 -356
rect -1366 -351 -1362 -350
rect -1725 -352 -1721 -351
rect -2092 -360 -2088 -359
rect -2059 -360 -2055 -359
rect -1818 -364 -1814 -363
rect -1333 -360 -1329 -359
rect -1333 -363 -1329 -362
rect -1818 -367 -1814 -366
rect -1366 -372 -1362 -371
rect -1366 -375 -1362 -374
rect -2092 -381 -2088 -380
rect -2092 -384 -2088 -383
rect -2059 -393 -2055 -392
rect -2059 -396 -2055 -395
rect -1366 -396 -1362 -395
rect -1366 -399 -1362 -398
rect -2092 -405 -2088 -404
rect -2092 -408 -2088 -407
rect -1366 -420 -1362 -419
rect -1333 -420 -1329 -419
rect -1366 -423 -1362 -422
rect -2092 -429 -2088 -428
rect -1333 -423 -1329 -422
rect -2092 -432 -2088 -431
rect -1366 -444 -1362 -443
rect -1366 -447 -1362 -446
rect -2092 -453 -2088 -452
rect -2059 -453 -2055 -452
rect -1544 -454 -1540 -453
rect -2092 -456 -2088 -455
rect -2059 -456 -2055 -455
rect -1485 -455 -1481 -450
rect -1544 -457 -1540 -456
rect -1485 -458 -1481 -457
rect -1366 -468 -1362 -467
rect -1349 -468 -1345 -467
rect -1333 -468 -1329 -467
rect -2092 -477 -2088 -476
rect -1825 -477 -1821 -476
rect -1792 -477 -1788 -476
rect -1366 -471 -1362 -470
rect -1349 -471 -1345 -470
rect -2092 -480 -2088 -479
rect -1825 -480 -1821 -479
rect -1792 -480 -1788 -479
rect -1333 -471 -1329 -470
rect -2092 -501 -2088 -500
rect -2075 -501 -2071 -500
rect -2059 -501 -2055 -500
rect -1825 -501 -1821 -500
rect -2092 -504 -2088 -503
rect -2075 -504 -2071 -503
rect -2059 -504 -2055 -503
rect -1825 -504 -1821 -503
rect -1792 -513 -1788 -512
rect -1638 -493 -1634 -492
rect -1621 -493 -1617 -492
rect -1638 -496 -1634 -495
rect -1621 -496 -1617 -495
rect -1541 -499 -1537 -498
rect -1519 -498 -1515 -497
rect -1273 -496 -1269 -495
rect -1273 -499 -1269 -498
rect -1541 -502 -1537 -501
rect -1519 -501 -1515 -500
rect -1792 -516 -1788 -515
rect -1999 -529 -1995 -528
rect -1825 -525 -1821 -524
rect -1620 -522 -1616 -521
rect -1620 -525 -1616 -524
rect -1825 -528 -1821 -527
rect -1999 -532 -1995 -531
rect -2092 -544 -2088 -543
rect -2092 -547 -2088 -546
rect -1825 -549 -1821 -548
rect -1825 -552 -1821 -551
rect -1366 -511 -1362 -510
rect -1366 -514 -1362 -513
rect -1519 -525 -1515 -524
rect -1541 -526 -1537 -525
rect -1541 -529 -1537 -528
rect -1519 -528 -1515 -527
rect -1825 -573 -1821 -572
rect -1792 -573 -1788 -572
rect -1825 -576 -1821 -575
rect -1792 -576 -1788 -575
rect -1825 -597 -1821 -596
rect -1825 -600 -1821 -599
rect -1825 -621 -1821 -620
rect -1808 -621 -1804 -620
rect -1792 -621 -1788 -620
rect -1825 -624 -1821 -623
rect -1808 -624 -1804 -623
rect -1792 -624 -1788 -623
rect -1732 -649 -1728 -648
rect -1732 -652 -1728 -651
rect -1825 -664 -1821 -663
rect -1825 -667 -1821 -666
<< pdiffusion >>
rect -2017 221 -2009 222
rect -1928 220 -1920 221
rect -2017 218 -2009 219
rect -2017 199 -2009 200
rect -2017 196 -2009 197
rect -1841 220 -1833 221
rect -1752 221 -1744 222
rect -1928 217 -1920 218
rect -1928 198 -1920 199
rect -1928 195 -1920 196
rect -1841 217 -1833 218
rect -1841 198 -1833 199
rect -1841 195 -1833 196
rect -1664 221 -1656 222
rect -1752 218 -1744 219
rect -1752 199 -1744 200
rect -1752 196 -1744 197
rect -1574 221 -1566 222
rect -1664 218 -1656 219
rect -1664 199 -1656 200
rect -1664 196 -1656 197
rect -1482 221 -1474 222
rect -1574 218 -1566 219
rect -1574 199 -1566 200
rect -1574 196 -1566 197
rect -1387 221 -1379 222
rect -1482 218 -1474 219
rect -1482 199 -1474 200
rect -1482 196 -1474 197
rect -1298 221 -1290 222
rect -1206 222 -1198 223
rect -1387 218 -1379 219
rect -1387 199 -1379 200
rect -1387 196 -1379 197
rect -1298 218 -1290 219
rect -1298 199 -1290 200
rect -1298 196 -1290 197
rect -1112 221 -1104 222
rect -1206 219 -1198 220
rect -1206 200 -1198 201
rect -1206 197 -1198 198
rect -1024 221 -1016 222
rect -1112 218 -1104 219
rect -1112 199 -1104 200
rect -1112 196 -1104 197
rect -934 221 -926 222
rect -1024 218 -1016 219
rect -1024 199 -1016 200
rect -1024 196 -1016 197
rect -843 221 -835 222
rect -934 218 -926 219
rect -934 199 -926 200
rect -934 196 -926 197
rect -752 221 -744 222
rect -843 218 -835 219
rect -843 199 -835 200
rect -843 196 -835 197
rect -663 221 -655 222
rect -752 218 -744 219
rect -752 199 -744 200
rect -752 196 -744 197
rect -663 218 -655 219
rect -663 199 -655 200
rect -663 196 -655 197
rect -2017 180 -2009 181
rect -1928 179 -1920 180
rect -1752 180 -1744 181
rect -1664 180 -1656 181
rect -1574 180 -1566 181
rect -1482 180 -1474 181
rect -1387 180 -1379 181
rect -1206 181 -1199 182
rect -1298 180 -1290 181
rect -1841 179 -1833 180
rect -2017 177 -2009 178
rect -1112 180 -1104 181
rect -1024 180 -1016 181
rect -934 180 -926 181
rect -843 180 -835 181
rect -752 180 -744 181
rect -663 180 -655 181
rect -1928 176 -1920 177
rect -1841 176 -1833 177
rect -1752 177 -1744 178
rect -1664 177 -1656 178
rect -1574 177 -1566 178
rect -1482 177 -1474 178
rect -1387 177 -1379 178
rect -1298 177 -1290 178
rect -1206 178 -1199 179
rect -1112 177 -1104 178
rect -1024 177 -1016 178
rect -934 177 -926 178
rect -843 177 -835 178
rect -752 177 -744 178
rect -663 177 -655 178
rect -1980 63 -1972 64
rect -826 66 -818 67
rect -767 65 -759 66
rect -1941 63 -1933 64
rect -1980 60 -1972 61
rect -1941 60 -1933 61
rect -826 63 -818 64
rect -767 62 -759 63
rect -1690 43 -1682 44
rect -1631 42 -1623 43
rect -1941 39 -1933 40
rect -1941 36 -1933 37
rect -1690 40 -1682 41
rect -1631 39 -1623 40
rect -899 39 -891 40
rect -1274 33 -1266 34
rect -1215 32 -1207 33
rect -1980 27 -1972 28
rect -1274 30 -1266 31
rect -1215 29 -1207 30
rect -1980 24 -1972 25
rect -1941 15 -1933 16
rect -1763 16 -1755 17
rect -1941 12 -1933 13
rect -2268 -15 -2260 -14
rect -1941 -9 -1933 -8
rect -2229 -15 -2221 -14
rect -1941 -12 -1933 -11
rect -1763 13 -1755 14
rect -899 36 -891 37
rect -794 22 -786 23
rect -768 22 -760 23
rect -899 17 -891 18
rect -899 14 -891 15
rect -1347 6 -1339 7
rect -1658 -1 -1650 0
rect -1632 -1 -1624 0
rect -1763 -6 -1755 -5
rect -1763 -9 -1755 -8
rect -2268 -18 -2260 -17
rect -2229 -18 -2221 -17
rect -1658 -4 -1650 -3
rect -1763 -25 -1755 -24
rect -1980 -33 -1972 -32
rect -1763 -28 -1755 -27
rect -1941 -33 -1933 -32
rect -2229 -39 -2221 -38
rect -2229 -42 -2221 -41
rect -1980 -36 -1972 -35
rect -1941 -36 -1933 -35
rect -2268 -51 -2260 -50
rect -2268 -54 -2260 -53
rect -1941 -57 -1933 -56
rect -2229 -63 -2221 -62
rect -1941 -60 -1933 -59
rect -2229 -66 -2221 -65
rect -1632 -4 -1624 -3
rect -794 19 -786 20
rect -1347 3 -1339 4
rect -899 -2 -891 -1
rect -1242 -11 -1234 -10
rect -899 -5 -891 -4
rect -1216 -11 -1208 -10
rect -1347 -16 -1339 -15
rect -1347 -19 -1339 -18
rect -1242 -14 -1234 -13
rect -1658 -35 -1650 -34
rect -1632 -35 -1624 -34
rect -1347 -35 -1339 -34
rect -1658 -38 -1650 -37
rect -1632 -38 -1624 -37
rect -1347 -38 -1339 -37
rect -1980 -81 -1972 -80
rect -1961 -81 -1953 -80
rect -1216 -14 -1208 -13
rect -1242 -45 -1234 -44
rect -1216 -45 -1208 -44
rect -768 19 -760 20
rect -794 -12 -786 -11
rect -768 -12 -760 -11
rect -794 -15 -786 -14
rect -768 -15 -760 -14
rect -1242 -48 -1234 -47
rect -1216 -48 -1208 -47
rect -1941 -81 -1933 -80
rect -2229 -87 -2221 -86
rect -2229 -90 -2221 -89
rect -1980 -84 -1972 -83
rect -1961 -84 -1953 -83
rect -1941 -84 -1933 -83
rect -1068 -88 -1060 -87
rect -1029 -88 -1021 -87
rect -1068 -91 -1060 -90
rect -1029 -91 -1021 -90
rect -2268 -111 -2260 -110
rect -1941 -109 -1933 -108
rect -2229 -111 -2221 -110
rect -2268 -114 -2260 -113
rect -2229 -114 -2221 -113
rect -1941 -112 -1933 -111
rect -1029 -112 -1021 -111
rect -1029 -115 -1021 -114
rect -2036 -124 -2028 -123
rect -2036 -127 -2028 -126
rect -1068 -124 -1060 -123
rect -2229 -135 -2221 -134
rect -1486 -137 -1478 -136
rect -1068 -127 -1060 -126
rect -1029 -136 -1021 -135
rect -1447 -137 -1439 -136
rect -2229 -138 -2221 -137
rect -1486 -140 -1478 -139
rect -1447 -140 -1439 -139
rect -1029 -139 -1021 -138
rect -2268 -159 -2260 -158
rect -2249 -159 -2241 -158
rect -2229 -159 -2221 -158
rect -1029 -160 -1021 -159
rect -1447 -161 -1439 -160
rect -2268 -162 -2260 -161
rect -2249 -162 -2241 -161
rect -2229 -162 -2221 -161
rect -1447 -164 -1439 -163
rect -1029 -163 -1021 -162
rect -1737 -177 -1729 -176
rect -1486 -173 -1478 -172
rect -1698 -177 -1690 -176
rect -1737 -180 -1729 -179
rect -1698 -180 -1690 -179
rect -1486 -176 -1478 -175
rect -1068 -184 -1060 -183
rect -1029 -184 -1021 -183
rect -1447 -185 -1439 -184
rect -2229 -187 -2221 -186
rect -2229 -190 -2221 -189
rect -1447 -188 -1439 -187
rect -1068 -187 -1060 -186
rect -1029 -187 -1021 -186
rect -1698 -201 -1690 -200
rect -2324 -202 -2316 -201
rect -2324 -205 -2316 -204
rect -1698 -204 -1690 -203
rect -1029 -208 -1021 -207
rect -1447 -209 -1439 -208
rect -1737 -213 -1729 -212
rect -1737 -216 -1729 -215
rect -1447 -212 -1439 -211
rect -1029 -211 -1021 -210
rect -1698 -225 -1690 -224
rect -1698 -228 -1690 -227
rect -1486 -233 -1478 -232
rect -1068 -232 -1060 -231
rect -1049 -232 -1041 -231
rect -1029 -232 -1021 -231
rect -1447 -233 -1439 -232
rect -1486 -236 -1478 -235
rect -1447 -236 -1439 -235
rect -1068 -235 -1060 -234
rect -1049 -235 -1041 -234
rect -1029 -235 -1021 -234
rect -1698 -249 -1690 -248
rect -1698 -252 -1690 -251
rect -1447 -257 -1439 -256
rect -1447 -260 -1439 -259
rect -1029 -260 -1021 -259
rect -1029 -263 -1021 -262
rect -1737 -273 -1729 -272
rect -1698 -273 -1690 -272
rect -1737 -276 -1729 -275
rect -1698 -276 -1690 -275
rect -1486 -281 -1478 -280
rect -1467 -281 -1459 -280
rect -1124 -275 -1116 -274
rect -1447 -281 -1439 -280
rect -1124 -278 -1116 -277
rect -1486 -284 -1478 -283
rect -1467 -284 -1459 -283
rect -1447 -284 -1439 -283
rect -1698 -297 -1690 -296
rect -1698 -300 -1690 -299
rect -1447 -309 -1439 -308
rect -1737 -321 -1729 -320
rect -1718 -321 -1710 -320
rect -1447 -312 -1439 -311
rect -1698 -321 -1690 -320
rect -1737 -324 -1729 -323
rect -1718 -324 -1710 -323
rect -1698 -324 -1690 -323
rect -1542 -324 -1534 -323
rect -1285 -324 -1277 -323
rect -1246 -324 -1238 -323
rect -1542 -327 -1534 -326
rect -1285 -327 -1277 -326
rect -1246 -327 -1238 -326
rect -1246 -348 -1238 -347
rect -1698 -349 -1690 -348
rect -2011 -357 -2003 -356
rect -1698 -352 -1690 -351
rect -1246 -351 -1238 -350
rect -1972 -357 -1964 -356
rect -2011 -360 -2003 -359
rect -1972 -360 -1964 -359
rect -1285 -360 -1277 -359
rect -1793 -364 -1785 -363
rect -1793 -367 -1785 -366
rect -1285 -363 -1277 -362
rect -1246 -372 -1238 -371
rect -1246 -375 -1238 -374
rect -1972 -381 -1964 -380
rect -1972 -384 -1964 -383
rect -2011 -393 -2003 -392
rect -2011 -396 -2003 -395
rect -1246 -396 -1238 -395
rect -1246 -399 -1238 -398
rect -1972 -405 -1964 -404
rect -1972 -408 -1964 -407
rect -1285 -420 -1277 -419
rect -1246 -420 -1238 -419
rect -1972 -429 -1964 -428
rect -1285 -423 -1277 -422
rect -1246 -423 -1238 -422
rect -1972 -432 -1964 -431
rect -1246 -444 -1238 -443
rect -2011 -453 -2003 -452
rect -1972 -453 -1964 -452
rect -1522 -454 -1514 -453
rect -2011 -456 -2003 -455
rect -1972 -456 -1964 -455
rect -1246 -447 -1238 -446
rect -1463 -455 -1455 -454
rect -1522 -457 -1514 -456
rect -1463 -458 -1455 -457
rect -1285 -468 -1277 -467
rect -1266 -468 -1258 -467
rect -1246 -468 -1238 -467
rect -1972 -477 -1964 -476
rect -1744 -477 -1736 -476
rect -1705 -477 -1697 -476
rect -1972 -480 -1964 -479
rect -1744 -480 -1736 -479
rect -1705 -480 -1697 -479
rect -1595 -481 -1587 -480
rect -1285 -471 -1277 -470
rect -1266 -471 -1258 -470
rect -1246 -471 -1238 -470
rect -2011 -501 -2003 -500
rect -1992 -501 -1984 -500
rect -1972 -501 -1964 -500
rect -1705 -501 -1697 -500
rect -2011 -504 -2003 -503
rect -1992 -504 -1984 -503
rect -1972 -504 -1964 -503
rect -1705 -504 -1697 -503
rect -1744 -513 -1736 -512
rect -1595 -484 -1587 -483
rect -1490 -498 -1482 -497
rect -1246 -496 -1238 -495
rect -1464 -498 -1456 -497
rect -1595 -503 -1587 -502
rect -1595 -506 -1587 -505
rect -1490 -501 -1482 -500
rect -1744 -516 -1736 -515
rect -1595 -522 -1587 -521
rect -1705 -525 -1697 -524
rect -1972 -529 -1964 -528
rect -1972 -532 -1964 -531
rect -1705 -528 -1697 -527
rect -1595 -525 -1587 -524
rect -2067 -544 -2059 -543
rect -2067 -547 -2059 -546
rect -1705 -549 -1697 -548
rect -1705 -552 -1697 -551
rect -1464 -501 -1456 -500
rect -1246 -499 -1238 -498
rect -1341 -511 -1333 -510
rect -1341 -514 -1333 -513
rect -1490 -532 -1482 -531
rect -1464 -532 -1456 -531
rect -1490 -535 -1482 -534
rect -1464 -535 -1456 -534
rect -1744 -573 -1736 -572
rect -1705 -573 -1697 -572
rect -1744 -576 -1736 -575
rect -1705 -576 -1697 -575
rect -1705 -597 -1697 -596
rect -1705 -600 -1697 -599
rect -1744 -621 -1736 -620
rect -1725 -621 -1717 -620
rect -1705 -621 -1697 -620
rect -1744 -624 -1736 -623
rect -1725 -624 -1717 -623
rect -1705 -624 -1697 -623
rect -1705 -649 -1697 -648
rect -1705 -652 -1697 -651
rect -1800 -664 -1792 -663
rect -1800 -667 -1792 -666
<< metal1 >>
rect -2056 226 -2052 250
rect -2031 225 -2027 250
rect -1967 225 -1963 249
rect -1942 224 -1938 249
rect -1880 225 -1876 249
rect -1855 224 -1851 249
rect -2028 214 -2017 218
rect -2050 210 -2043 214
rect -2050 206 -2047 210
rect -2028 206 -2024 214
rect -1939 213 -1928 217
rect -1852 213 -1841 217
rect -1961 209 -1954 213
rect -2056 202 -2047 206
rect -2039 202 -2024 206
rect -1961 205 -1958 209
rect -1939 205 -1935 213
rect -1874 209 -1867 213
rect -1874 205 -1871 209
rect -1852 205 -1848 213
rect -2028 196 -2024 202
rect -1967 201 -1958 205
rect -1950 201 -1935 205
rect -2028 192 -2017 196
rect -1939 195 -1935 201
rect -1880 201 -1871 205
rect -1863 201 -1848 205
rect -1852 195 -1848 201
rect -2028 184 -2024 192
rect -1939 191 -1928 195
rect -1852 191 -1841 195
rect -1939 183 -1935 191
rect -1852 183 -1848 191
rect -2038 173 -2017 177
rect -2030 154 -2026 173
rect -1949 172 -1928 176
rect -1862 172 -1841 176
rect -2332 150 -2026 154
rect -2332 37 -2328 150
rect -1941 124 -1937 172
rect -2044 120 -1937 124
rect -2288 49 -2086 53
rect -2288 37 -2284 49
rect -2332 -27 -2328 33
rect -2288 12 -2284 33
rect -2243 12 -2183 16
rect -2288 8 -2276 12
rect -2288 -11 -2284 8
rect -2332 -31 -2298 -27
rect -2332 -75 -2328 -31
rect -2302 -47 -2298 -31
rect -2280 -33 -2276 8
rect -2250 8 -2239 12
rect -2250 -26 -2246 8
rect -2243 -1 -2239 8
rect -2250 -30 -2235 -26
rect -2280 -37 -2253 -33
rect -2280 -59 -2276 -37
rect -2332 -83 -2328 -79
rect -2257 -98 -2253 -37
rect -2250 -35 -2246 -30
rect -2239 -98 -2235 -30
rect -2340 -102 -2300 -98
rect -2340 -198 -2336 -102
rect -2304 -107 -2300 -102
rect -2257 -102 -2246 -98
rect -2312 -118 -2268 -114
rect -2294 -162 -2290 -118
rect -2257 -131 -2253 -102
rect -2250 -145 -2246 -102
rect -2239 -102 -2210 -98
rect -2239 -107 -2235 -102
rect -2312 -166 -2268 -162
rect -2294 -176 -2290 -166
rect -2214 -169 -2210 -102
rect -2246 -173 -2210 -169
rect -2294 -179 -2241 -176
rect -2245 -183 -2241 -179
rect -2252 -194 -2229 -190
rect -2345 -209 -2324 -205
rect -2339 -234 -2334 -209
rect -2245 -226 -2241 -194
rect -2187 -571 -2183 12
rect -2090 -140 -2086 49
rect -2044 51 -2040 120
rect -1854 111 -1850 172
rect -2000 107 -1850 111
rect -2000 90 -1996 107
rect -1955 90 -1853 94
rect -2000 86 -1988 90
rect -2000 67 -1996 86
rect -2044 47 -2010 51
rect -2044 3 -2040 47
rect -2014 31 -2010 47
rect -1992 45 -1988 86
rect -1962 86 -1951 90
rect -1962 52 -1958 86
rect -1955 77 -1951 86
rect -1962 48 -1947 52
rect -1992 41 -1965 45
rect -1992 19 -1988 41
rect -2044 -5 -2040 -1
rect -1969 -20 -1965 41
rect -1962 43 -1958 48
rect -1951 -20 -1947 48
rect -2052 -24 -2012 -20
rect -2052 -120 -2048 -24
rect -2016 -29 -2012 -24
rect -1969 -24 -1958 -20
rect -2024 -40 -1980 -36
rect -2006 -84 -2002 -40
rect -1969 -53 -1965 -24
rect -1962 -67 -1958 -24
rect -1951 -24 -1922 -20
rect -1951 -29 -1947 -24
rect -2024 -88 -1980 -84
rect -2006 -98 -2002 -88
rect -1926 -91 -1922 -24
rect -1958 -95 -1922 -91
rect -2006 -101 -1953 -98
rect -1957 -105 -1953 -101
rect -1964 -116 -1941 -112
rect -2057 -131 -2036 -127
rect -2051 -140 -2046 -131
rect -2090 -144 -2046 -140
rect -1957 -199 -1953 -116
rect -2075 -203 -1953 -199
rect -2075 -369 -2071 -203
rect -2031 -293 -1866 -289
rect -2031 -330 -2027 -293
rect -1986 -330 -1894 -326
rect -2031 -334 -2019 -330
rect -2031 -353 -2027 -334
rect -2075 -373 -2041 -369
rect -2075 -417 -2071 -373
rect -2045 -389 -2041 -373
rect -2023 -375 -2019 -334
rect -1993 -334 -1982 -330
rect -1993 -368 -1989 -334
rect -1986 -343 -1982 -334
rect -1993 -372 -1978 -368
rect -2023 -379 -1996 -375
rect -2023 -401 -2019 -379
rect -2075 -425 -2071 -421
rect -2000 -440 -1996 -379
rect -1993 -377 -1989 -372
rect -1982 -440 -1978 -372
rect -2083 -444 -2043 -440
rect -2083 -540 -2079 -444
rect -2047 -449 -2043 -444
rect -2000 -444 -1989 -440
rect -2055 -460 -2011 -456
rect -2037 -504 -2033 -460
rect -2000 -473 -1996 -444
rect -1993 -487 -1989 -444
rect -1982 -444 -1953 -440
rect -1982 -449 -1978 -444
rect -2055 -508 -2011 -504
rect -2037 -518 -2033 -508
rect -1957 -511 -1953 -444
rect -1989 -515 -1953 -511
rect -2037 -521 -1984 -518
rect -1988 -525 -1984 -521
rect -1995 -536 -1972 -532
rect -2088 -551 -2067 -547
rect -2082 -571 -2077 -551
rect -2187 -576 -2076 -571
rect -1988 -729 -1984 -536
rect -1898 -705 -1894 -330
rect -1870 -692 -1866 -293
rect -1857 -392 -1853 90
rect -1838 -113 -1834 109
rect -1828 -105 -1824 133
rect -1814 9 -1810 242
rect -1791 226 -1787 250
rect -1766 225 -1762 250
rect -1703 226 -1699 250
rect -1678 225 -1674 250
rect -1613 226 -1609 250
rect -1588 225 -1584 250
rect -1521 226 -1517 250
rect -1496 225 -1492 250
rect -1426 226 -1422 250
rect -1401 225 -1397 250
rect -1763 214 -1752 218
rect -1675 214 -1664 218
rect -1585 214 -1574 218
rect -1493 214 -1482 218
rect -1398 214 -1387 218
rect -1785 210 -1778 214
rect -1785 206 -1782 210
rect -1763 206 -1759 214
rect -1697 210 -1690 214
rect -1697 206 -1694 210
rect -1675 206 -1671 214
rect -1607 210 -1600 214
rect -1607 206 -1604 210
rect -1585 206 -1581 214
rect -1515 210 -1508 214
rect -1515 206 -1512 210
rect -1493 206 -1489 214
rect -1420 210 -1413 214
rect -1420 206 -1417 210
rect -1398 206 -1394 214
rect -1791 202 -1782 206
rect -1774 202 -1759 206
rect -1763 196 -1759 202
rect -1703 202 -1694 206
rect -1686 202 -1671 206
rect -1675 196 -1671 202
rect -1613 202 -1604 206
rect -1596 202 -1581 206
rect -1585 196 -1581 202
rect -1521 202 -1512 206
rect -1504 202 -1489 206
rect -1493 196 -1489 202
rect -1426 202 -1417 206
rect -1409 202 -1394 206
rect -1398 196 -1394 202
rect -1763 192 -1752 196
rect -1675 192 -1664 196
rect -1585 192 -1574 196
rect -1493 192 -1482 196
rect -1398 192 -1387 196
rect -1763 184 -1759 192
rect -1675 184 -1671 192
rect -1585 184 -1581 192
rect -1493 184 -1489 192
rect -1398 184 -1394 192
rect -1773 173 -1752 177
rect -1685 173 -1664 177
rect -1595 173 -1574 177
rect -1503 173 -1482 177
rect -1408 173 -1387 177
rect -1765 152 -1761 173
rect -1677 137 -1673 173
rect -1587 160 -1583 173
rect -1628 156 -1583 160
rect -1628 127 -1624 156
rect -1495 150 -1491 173
rect -1765 123 -1624 127
rect -1587 146 -1491 150
rect -1765 113 -1761 123
rect -1587 115 -1583 146
rect -1400 141 -1396 173
rect -1362 154 -1358 242
rect -1337 226 -1333 250
rect -1312 225 -1308 250
rect -1245 227 -1241 251
rect -1220 226 -1216 251
rect -1151 226 -1147 250
rect -1126 225 -1122 250
rect -1063 226 -1059 250
rect -1038 225 -1034 250
rect -973 226 -969 250
rect -948 225 -944 250
rect -1309 214 -1298 218
rect -1217 215 -1206 219
rect -1331 210 -1324 214
rect -1331 206 -1328 210
rect -1309 206 -1305 214
rect -1239 211 -1232 215
rect -1239 207 -1236 211
rect -1217 207 -1213 215
rect -1123 214 -1112 218
rect -1035 214 -1024 218
rect -945 214 -934 218
rect -1145 210 -1138 214
rect -1337 202 -1328 206
rect -1320 202 -1305 206
rect -1309 196 -1305 202
rect -1245 203 -1236 207
rect -1228 203 -1213 207
rect -1145 206 -1142 210
rect -1123 206 -1119 214
rect -1057 210 -1050 214
rect -1057 206 -1054 210
rect -1035 206 -1031 214
rect -967 210 -960 214
rect -967 206 -964 210
rect -945 206 -941 214
rect -1217 197 -1213 203
rect -1151 202 -1142 206
rect -1134 202 -1119 206
rect -1309 192 -1298 196
rect -1217 193 -1206 197
rect -1123 196 -1119 202
rect -1063 202 -1054 206
rect -1046 202 -1031 206
rect -1035 196 -1031 202
rect -973 202 -964 206
rect -956 202 -941 206
rect -945 196 -941 202
rect -1309 184 -1305 192
rect -1217 185 -1213 193
rect -1123 192 -1112 196
rect -1035 192 -1024 196
rect -945 192 -934 196
rect -1123 184 -1119 192
rect -1035 184 -1031 192
rect -945 184 -941 192
rect -1319 173 -1298 177
rect -1227 174 -1206 178
rect -1777 109 -1761 113
rect -1703 111 -1583 115
rect -1558 137 -1396 141
rect -1802 21 -1798 94
rect -1703 82 -1699 111
rect -1558 107 -1554 137
rect -1311 131 -1307 173
rect -1414 127 -1307 131
rect -1219 121 -1215 174
rect -1133 173 -1112 177
rect -1045 173 -1024 177
rect -955 173 -934 177
rect -1777 77 -1699 82
rect -1777 20 -1773 77
rect -1703 61 -1699 77
rect -1727 58 -1720 61
rect -1716 58 -1699 61
rect -1727 14 -1724 58
rect -1703 47 -1699 58
rect -1644 103 -1554 107
rect -1506 117 -1215 121
rect -1644 98 -1640 103
rect -1644 67 -1640 94
rect -1644 63 -1602 67
rect -1644 46 -1640 63
rect -1774 9 -1763 13
rect -1727 10 -1705 14
rect -1796 5 -1789 9
rect -1796 1 -1793 5
rect -1774 1 -1770 9
rect -1802 -3 -1793 1
rect -1785 -3 -1770 1
rect -1696 0 -1687 4
rect -1650 0 -1639 4
rect -1774 -9 -1770 -3
rect -1696 -5 -1693 0
rect -1642 -4 -1639 0
rect -1705 -9 -1693 -5
rect -1683 -8 -1658 -4
rect -1642 -8 -1632 -4
rect -1774 -13 -1763 -9
rect -1774 -21 -1770 -13
rect -1696 -27 -1687 -23
rect -1784 -32 -1763 -28
rect -1696 -32 -1693 -27
rect -1678 -31 -1673 -8
rect -1776 -86 -1772 -32
rect -1705 -36 -1693 -32
rect -1683 -35 -1673 -31
rect -1650 -34 -1638 -30
rect -1747 -78 -1741 -39
rect -1678 -38 -1673 -35
rect -1641 -38 -1638 -34
rect -1678 -42 -1658 -38
rect -1641 -42 -1632 -38
rect -1776 -91 -1708 -86
rect -1828 -109 -1753 -105
rect -1838 -116 -1797 -113
rect -1801 -189 -1797 -116
rect -1757 -150 -1753 -109
rect -1712 -150 -1708 -91
rect -1678 -103 -1673 -42
rect -1607 -60 -1602 63
rect -1630 -64 -1602 -60
rect -1588 -76 -1546 -73
rect -1588 -103 -1584 -76
rect -1550 -85 -1546 -76
rect -1506 -85 -1502 117
rect -1287 100 -1141 104
rect -1398 -1 -1394 80
rect -1386 11 -1382 84
rect -1287 72 -1283 100
rect -1125 93 -1121 173
rect -1037 104 -1033 173
rect -947 155 -943 173
rect -1062 100 -1033 104
rect -991 151 -943 155
rect -991 96 -987 151
rect -907 148 -903 242
rect -882 226 -878 250
rect -857 225 -853 250
rect -791 226 -787 250
rect -766 225 -762 250
rect -702 226 -698 250
rect -677 225 -673 250
rect -854 214 -843 218
rect -763 214 -752 218
rect -674 214 -663 218
rect -876 210 -869 214
rect -876 206 -873 210
rect -854 206 -850 214
rect -785 210 -778 214
rect -785 206 -782 210
rect -763 206 -759 214
rect -696 210 -689 214
rect -696 206 -693 210
rect -674 206 -670 214
rect -882 202 -873 206
rect -865 202 -850 206
rect -854 196 -850 202
rect -791 202 -782 206
rect -774 202 -759 206
rect -763 196 -759 202
rect -702 202 -693 206
rect -685 202 -670 206
rect -674 196 -670 202
rect -854 192 -843 196
rect -763 192 -752 196
rect -674 192 -663 196
rect -854 184 -850 192
rect -763 184 -759 192
rect -674 184 -670 192
rect -864 173 -843 177
rect -773 173 -752 177
rect -684 173 -663 177
rect -1361 67 -1283 72
rect -1361 10 -1357 67
rect -1287 51 -1283 67
rect -1311 48 -1304 51
rect -1300 48 -1283 51
rect -1311 4 -1308 48
rect -1287 37 -1283 48
rect -1228 89 -1121 93
rect -1088 92 -987 96
rect -950 144 -903 148
rect -856 151 -852 173
rect -856 147 -835 151
rect -765 149 -761 173
rect -1228 88 -1224 89
rect -1228 57 -1224 84
rect -1228 53 -1186 57
rect -1228 36 -1224 53
rect -1358 -1 -1347 3
rect -1311 0 -1289 4
rect -1380 -5 -1373 -1
rect -1380 -9 -1377 -5
rect -1358 -9 -1354 -1
rect -1386 -13 -1377 -9
rect -1369 -13 -1354 -9
rect -1280 -10 -1271 -6
rect -1234 -10 -1223 -6
rect -1358 -19 -1354 -13
rect -1280 -15 -1277 -10
rect -1226 -14 -1223 -10
rect -1289 -19 -1277 -15
rect -1267 -18 -1242 -14
rect -1226 -18 -1216 -14
rect -1358 -23 -1347 -19
rect -1358 -31 -1354 -23
rect -1280 -37 -1271 -33
rect -1368 -42 -1347 -38
rect -1280 -42 -1277 -37
rect -1262 -41 -1257 -18
rect -1678 -107 -1584 -103
rect -1757 -154 -1745 -150
rect -1757 -173 -1753 -154
rect -1801 -193 -1767 -189
rect -1801 -237 -1797 -193
rect -1771 -209 -1767 -193
rect -1749 -195 -1745 -154
rect -1719 -154 -1708 -150
rect -1719 -188 -1715 -154
rect -1712 -163 -1708 -154
rect -1550 -149 -1546 -89
rect -1506 -110 -1502 -89
rect -1419 -94 -1414 -81
rect -1360 -106 -1356 -42
rect -1289 -46 -1277 -42
rect -1267 -45 -1257 -41
rect -1234 -44 -1222 -40
rect -1331 -88 -1325 -49
rect -1262 -48 -1257 -45
rect -1225 -48 -1222 -44
rect -1262 -52 -1242 -48
rect -1225 -52 -1216 -48
rect -1461 -110 -1356 -106
rect -1506 -114 -1494 -110
rect -1506 -133 -1502 -114
rect -1550 -153 -1516 -149
rect -1719 -192 -1704 -188
rect -1749 -199 -1722 -195
rect -1749 -221 -1745 -199
rect -1801 -245 -1797 -241
rect -1726 -260 -1722 -199
rect -1719 -197 -1715 -192
rect -1708 -260 -1704 -192
rect -1550 -197 -1546 -153
rect -1520 -169 -1516 -153
rect -1498 -155 -1494 -114
rect -1468 -114 -1457 -110
rect -1468 -148 -1464 -114
rect -1461 -123 -1457 -114
rect -1419 -136 -1414 -118
rect -1262 -120 -1257 -52
rect -1191 -70 -1186 53
rect -1214 -74 -1186 -70
rect -1175 -27 -1128 -24
rect -1175 -120 -1171 -27
rect -1132 -36 -1128 -27
rect -1088 -36 -1084 92
rect -950 32 -946 144
rect -938 44 -934 117
rect -839 105 -835 147
rect -913 100 -835 105
rect -913 43 -909 100
rect -839 84 -835 100
rect -863 81 -856 84
rect -852 81 -835 84
rect -863 37 -860 81
rect -839 70 -835 81
rect -780 145 -761 149
rect -780 121 -776 145
rect -780 90 -776 117
rect -780 86 -738 90
rect -780 69 -776 86
rect -910 32 -899 36
rect -863 33 -841 37
rect -932 28 -925 32
rect -932 24 -929 28
rect -910 24 -906 32
rect -938 20 -929 24
rect -921 20 -906 24
rect -832 23 -823 27
rect -786 23 -775 27
rect -910 14 -906 20
rect -832 18 -829 23
rect -778 19 -775 23
rect -841 14 -829 18
rect -819 15 -794 19
rect -778 15 -768 19
rect -910 10 -899 14
rect -910 2 -906 10
rect -832 -4 -823 0
rect -920 -9 -899 -5
rect -832 -9 -829 -4
rect -814 -8 -809 15
rect -1132 -100 -1128 -40
rect -1088 -61 -1084 -40
rect -912 -57 -908 -9
rect -1043 -61 -908 -57
rect -841 -13 -829 -9
rect -819 -12 -809 -8
rect -786 -11 -774 -7
rect -883 -55 -877 -16
rect -814 -15 -809 -12
rect -777 -15 -774 -11
rect -814 -19 -794 -15
rect -777 -19 -768 -15
rect -1088 -65 -1076 -61
rect -1088 -84 -1084 -65
rect -1132 -104 -1098 -100
rect -1262 -123 -1171 -120
rect -1419 -140 -1301 -136
rect -1468 -152 -1453 -148
rect -1498 -159 -1471 -155
rect -1498 -181 -1494 -159
rect -1550 -205 -1546 -201
rect -1475 -220 -1471 -159
rect -1468 -157 -1464 -152
rect -1457 -220 -1453 -152
rect -1558 -224 -1518 -220
rect -1809 -264 -1769 -260
rect -1809 -360 -1805 -264
rect -1773 -269 -1769 -264
rect -1726 -264 -1715 -260
rect -1781 -280 -1737 -276
rect -1763 -324 -1759 -280
rect -1726 -293 -1722 -264
rect -1719 -307 -1715 -264
rect -1708 -264 -1679 -260
rect -1708 -269 -1704 -264
rect -1781 -328 -1737 -324
rect -1763 -338 -1759 -328
rect -1683 -331 -1679 -264
rect -1715 -335 -1679 -331
rect -1646 -323 -1578 -319
rect -1558 -320 -1554 -224
rect -1522 -229 -1518 -224
rect -1475 -224 -1464 -220
rect -1530 -240 -1486 -236
rect -1512 -284 -1508 -240
rect -1475 -253 -1471 -224
rect -1468 -267 -1464 -224
rect -1457 -224 -1428 -220
rect -1457 -229 -1453 -224
rect -1530 -288 -1486 -284
rect -1512 -298 -1508 -288
rect -1432 -291 -1428 -224
rect -1464 -295 -1428 -291
rect -1393 -263 -1345 -260
rect -1512 -301 -1459 -298
rect -1463 -305 -1459 -301
rect -1470 -316 -1447 -312
rect -1763 -341 -1710 -338
rect -1714 -345 -1710 -341
rect -1721 -356 -1698 -352
rect -1814 -371 -1793 -367
rect -1808 -392 -1803 -371
rect -1714 -383 -1710 -356
rect -1857 -396 -1803 -392
rect -1764 -387 -1710 -383
rect -1844 -417 -1804 -413
rect -1808 -489 -1804 -417
rect -1764 -450 -1760 -387
rect -1719 -450 -1664 -446
rect -1764 -454 -1752 -450
rect -1764 -473 -1760 -454
rect -1808 -493 -1774 -489
rect -1808 -537 -1804 -493
rect -1778 -509 -1774 -493
rect -1756 -495 -1752 -454
rect -1726 -454 -1715 -450
rect -1726 -488 -1722 -454
rect -1719 -463 -1715 -454
rect -1646 -488 -1642 -323
rect -1563 -331 -1542 -327
rect -1557 -351 -1552 -331
rect -1463 -344 -1459 -316
rect -1393 -344 -1389 -263
rect -1349 -272 -1345 -263
rect -1305 -272 -1301 -140
rect -1132 -148 -1128 -104
rect -1102 -120 -1098 -104
rect -1080 -106 -1076 -65
rect -1050 -65 -1039 -61
rect -1050 -99 -1046 -65
rect -1043 -74 -1039 -65
rect -1050 -103 -1035 -99
rect -1080 -110 -1053 -106
rect -1080 -132 -1076 -110
rect -1132 -156 -1128 -152
rect -1057 -171 -1053 -110
rect -1050 -108 -1046 -103
rect -1039 -171 -1035 -103
rect -1140 -175 -1100 -171
rect -1140 -271 -1136 -175
rect -1104 -180 -1100 -175
rect -1057 -175 -1046 -171
rect -1112 -191 -1068 -187
rect -1094 -235 -1090 -191
rect -1057 -204 -1053 -175
rect -1050 -218 -1046 -175
rect -1039 -175 -1010 -171
rect -1039 -180 -1035 -175
rect -1112 -239 -1068 -235
rect -1094 -249 -1090 -239
rect -1014 -242 -1010 -175
rect -1046 -246 -1010 -242
rect -1094 -252 -1041 -249
rect -1045 -256 -1041 -252
rect -1052 -267 -1029 -263
rect -1349 -336 -1345 -276
rect -1305 -297 -1301 -276
rect -1145 -282 -1124 -278
rect -1139 -293 -1134 -282
rect -1260 -297 -1134 -293
rect -1305 -301 -1293 -297
rect -1305 -320 -1301 -301
rect -1349 -340 -1315 -336
rect -1463 -348 -1389 -344
rect -1349 -384 -1345 -340
rect -1319 -356 -1315 -340
rect -1297 -342 -1293 -301
rect -1267 -301 -1256 -297
rect -1267 -335 -1263 -301
rect -1260 -310 -1256 -301
rect -1267 -339 -1252 -335
rect -1297 -346 -1270 -342
rect -1297 -368 -1293 -346
rect -1634 -476 -1630 -403
rect -1535 -415 -1531 -394
rect -1609 -420 -1531 -415
rect -1609 -477 -1605 -420
rect -1535 -436 -1531 -420
rect -1559 -439 -1552 -436
rect -1548 -439 -1531 -436
rect -1559 -483 -1556 -439
rect -1535 -450 -1531 -439
rect -1476 -394 -1395 -390
rect -1476 -399 -1472 -394
rect -1476 -430 -1472 -403
rect -1476 -434 -1434 -430
rect -1476 -451 -1472 -434
rect -1606 -488 -1595 -484
rect -1559 -487 -1537 -483
rect -1726 -492 -1711 -488
rect -1628 -492 -1621 -488
rect -1756 -499 -1729 -495
rect -1756 -521 -1752 -499
rect -1808 -545 -1804 -541
rect -1733 -560 -1729 -499
rect -1726 -497 -1722 -492
rect -1715 -560 -1711 -492
rect -1628 -496 -1625 -492
rect -1606 -496 -1602 -488
rect -1634 -500 -1625 -496
rect -1617 -500 -1602 -496
rect -1528 -497 -1519 -493
rect -1482 -497 -1471 -493
rect -1606 -506 -1602 -500
rect -1528 -502 -1525 -497
rect -1474 -501 -1471 -497
rect -1537 -506 -1525 -502
rect -1515 -505 -1490 -501
rect -1474 -505 -1464 -501
rect -1606 -510 -1595 -506
rect -1606 -518 -1602 -510
rect -1528 -524 -1519 -520
rect -1616 -529 -1595 -525
rect -1528 -529 -1525 -524
rect -1510 -528 -1505 -505
rect -1816 -564 -1776 -560
rect -1816 -660 -1812 -564
rect -1780 -569 -1776 -564
rect -1733 -564 -1722 -560
rect -1788 -580 -1744 -576
rect -1770 -624 -1766 -580
rect -1733 -593 -1729 -564
rect -1726 -607 -1722 -564
rect -1715 -564 -1686 -560
rect -1715 -569 -1711 -564
rect -1788 -628 -1744 -624
rect -1770 -638 -1766 -628
rect -1690 -631 -1686 -564
rect -1608 -577 -1604 -529
rect -1722 -635 -1686 -631
rect -1654 -581 -1604 -577
rect -1537 -533 -1525 -529
rect -1515 -532 -1505 -528
rect -1482 -531 -1470 -527
rect -1579 -575 -1573 -536
rect -1510 -535 -1505 -532
rect -1473 -535 -1470 -531
rect -1510 -539 -1490 -535
rect -1473 -539 -1464 -535
rect -1770 -641 -1717 -638
rect -1721 -645 -1717 -641
rect -1728 -656 -1705 -652
rect -1821 -671 -1800 -667
rect -1815 -692 -1810 -671
rect -1721 -684 -1717 -656
rect -1870 -696 -1810 -692
rect -1654 -705 -1650 -581
rect -1510 -640 -1505 -539
rect -1439 -557 -1434 -434
rect -1399 -539 -1395 -394
rect -1349 -392 -1345 -388
rect -1274 -407 -1270 -346
rect -1267 -344 -1263 -339
rect -1256 -407 -1252 -339
rect -1357 -411 -1317 -407
rect -1357 -507 -1353 -411
rect -1321 -416 -1317 -411
rect -1274 -411 -1263 -407
rect -1329 -427 -1285 -423
rect -1311 -471 -1307 -427
rect -1274 -440 -1270 -411
rect -1267 -454 -1263 -411
rect -1256 -411 -1227 -407
rect -1256 -416 -1252 -411
rect -1329 -475 -1285 -471
rect -1311 -485 -1307 -475
rect -1231 -478 -1227 -411
rect -1263 -482 -1227 -478
rect -1311 -488 -1258 -485
rect -1262 -492 -1258 -488
rect -1269 -503 -1246 -499
rect -1362 -518 -1341 -514
rect -1356 -539 -1351 -518
rect -1399 -543 -1351 -539
rect -1462 -561 -1434 -557
rect -1262 -635 -1258 -503
rect -1045 -560 -1041 -267
rect -814 -570 -809 -19
rect -743 -37 -738 86
rect -766 -41 -738 -37
rect -676 -570 -672 173
rect -1898 -709 -1650 -705
<< metal2 >>
rect -2068 242 -1814 246
rect -1810 242 -1362 246
rect -1358 242 -907 246
rect -903 242 -710 246
rect -2068 214 -2064 242
rect -2001 226 -1995 237
rect -2017 222 -1995 226
rect -2068 210 -2056 214
rect -2068 185 -2064 210
rect -2001 204 -1995 222
rect -2017 200 -1995 204
rect -2001 185 -1995 200
rect -2072 181 -2038 185
rect -2017 181 -1995 185
rect -2072 68 -2068 181
rect -2001 166 -1995 181
rect -1979 213 -1975 242
rect -1912 225 -1906 236
rect -1928 221 -1906 225
rect -1979 209 -1967 213
rect -1979 184 -1975 209
rect -1912 203 -1906 221
rect -1928 199 -1906 203
rect -1912 184 -1906 199
rect -1979 180 -1949 184
rect -1928 180 -1906 184
rect -1892 213 -1888 242
rect -1825 225 -1819 236
rect -1841 221 -1819 225
rect -1892 209 -1880 213
rect -1892 184 -1888 209
rect -1825 203 -1819 221
rect -1841 199 -1819 203
rect -1825 184 -1819 199
rect -1892 180 -1862 184
rect -1841 180 -1819 184
rect -1803 214 -1799 242
rect -1736 226 -1730 237
rect -1752 222 -1730 226
rect -1803 210 -1791 214
rect -1803 185 -1799 210
rect -1736 204 -1730 222
rect -1752 200 -1730 204
rect -1736 185 -1730 200
rect -1803 181 -1773 185
rect -1752 181 -1730 185
rect -1715 214 -1711 242
rect -1648 226 -1642 237
rect -1664 222 -1642 226
rect -1715 210 -1703 214
rect -1715 185 -1711 210
rect -1648 204 -1642 222
rect -1664 200 -1642 204
rect -1648 185 -1642 200
rect -1715 181 -1685 185
rect -1664 181 -1642 185
rect -1625 214 -1621 242
rect -1558 226 -1552 237
rect -1574 222 -1552 226
rect -1625 210 -1613 214
rect -1625 185 -1621 210
rect -1558 204 -1552 222
rect -1574 200 -1552 204
rect -1558 185 -1552 200
rect -1625 181 -1595 185
rect -1574 181 -1552 185
rect -1533 214 -1529 242
rect -1466 226 -1460 237
rect -1482 222 -1460 226
rect -1533 210 -1521 214
rect -1533 185 -1529 210
rect -1466 204 -1460 222
rect -1482 200 -1460 204
rect -1466 185 -1460 200
rect -1533 181 -1503 185
rect -1482 181 -1460 185
rect -1438 214 -1434 242
rect -1371 226 -1365 237
rect -1387 222 -1365 226
rect -1438 210 -1426 214
rect -1438 185 -1434 210
rect -1371 204 -1365 222
rect -1387 200 -1365 204
rect -1371 185 -1365 200
rect -1438 181 -1408 185
rect -1387 181 -1365 185
rect -1349 214 -1345 242
rect -1282 226 -1276 237
rect -1298 222 -1276 226
rect -1349 210 -1337 214
rect -1349 185 -1345 210
rect -1282 204 -1276 222
rect -1298 200 -1276 204
rect -1282 185 -1276 200
rect -1349 181 -1319 185
rect -1298 181 -1276 185
rect -1257 215 -1253 242
rect -1190 227 -1184 238
rect -1206 223 -1184 227
rect -1257 211 -1245 215
rect -1257 186 -1253 211
rect -1190 205 -1184 223
rect -1206 201 -1184 205
rect -1190 186 -1184 201
rect -1257 182 -1227 186
rect -1206 182 -1184 186
rect -2000 163 -1995 166
rect -1912 163 -1906 180
rect -1825 163 -1819 180
rect -1736 163 -1730 181
rect -1648 163 -1642 181
rect -1558 163 -1552 181
rect -1466 163 -1460 181
rect -1371 163 -1365 181
rect -1282 163 -1276 181
rect -1190 163 -1184 182
rect -1163 214 -1159 242
rect -1096 226 -1090 237
rect -1112 222 -1090 226
rect -1163 210 -1151 214
rect -1163 185 -1159 210
rect -1096 204 -1090 222
rect -1112 200 -1090 204
rect -1096 185 -1090 200
rect -1163 181 -1133 185
rect -1112 181 -1090 185
rect -1075 214 -1071 242
rect -1008 226 -1002 237
rect -1024 222 -1002 226
rect -1075 210 -1063 214
rect -1075 185 -1071 210
rect -1008 204 -1002 222
rect -1024 200 -1002 204
rect -1008 185 -1002 200
rect -1075 181 -1045 185
rect -1024 181 -1002 185
rect -985 214 -981 242
rect -918 226 -912 237
rect -934 222 -912 226
rect -985 210 -973 214
rect -985 185 -981 210
rect -918 204 -912 222
rect -934 200 -912 204
rect -918 185 -912 200
rect -985 181 -955 185
rect -934 181 -912 185
rect -894 214 -890 242
rect -827 226 -821 237
rect -843 222 -821 226
rect -894 210 -882 214
rect -894 185 -890 210
rect -827 204 -821 222
rect -843 200 -821 204
rect -827 185 -821 200
rect -894 181 -864 185
rect -843 181 -821 185
rect -803 214 -799 242
rect -736 226 -730 237
rect -752 222 -730 226
rect -803 210 -791 214
rect -803 185 -799 210
rect -736 204 -730 222
rect -752 200 -730 204
rect -736 185 -730 200
rect -803 181 -773 185
rect -752 181 -730 185
rect -714 214 -710 242
rect -647 226 -641 237
rect -663 222 -641 226
rect -714 210 -702 214
rect -714 185 -710 210
rect -647 204 -641 222
rect -663 200 -641 204
rect -647 185 -641 200
rect -714 181 -684 185
rect -663 181 -641 185
rect -1096 163 -1090 181
rect -1008 163 -1002 181
rect -918 163 -912 181
rect -827 163 -821 181
rect -736 163 -730 181
rect -647 163 -641 181
rect -2000 159 -641 163
rect -1922 74 -1918 159
rect -1928 68 -1918 74
rect -2072 64 -2057 68
rect -2043 64 -2024 68
rect -1980 64 -1954 68
rect -1941 64 -1918 68
rect -2072 44 -2068 64
rect -2043 60 -2040 64
rect -1957 60 -1954 64
rect -2061 56 -2040 60
rect -2028 56 -1972 60
rect -1957 56 -1933 60
rect -2072 40 -2057 44
rect -2072 37 -2068 40
rect -2360 33 -2068 37
rect -2360 -10 -2356 33
rect -2072 20 -2068 33
rect -2061 32 -2040 36
rect -2043 28 -2024 32
rect -2072 16 -2057 20
rect -2072 -4 -2068 16
rect -2043 12 -2040 28
rect -2006 24 -2002 56
rect -1928 44 -1918 64
rect -1941 40 -1918 44
rect -1957 32 -1933 36
rect -1980 28 -1954 32
rect -2028 20 -1972 24
rect -2061 8 -2040 12
rect -2040 -1 -2016 3
rect -2216 -8 -2126 -4
rect -2216 -10 -2206 -8
rect -2360 -14 -2345 -10
rect -2331 -14 -2312 -10
rect -2268 -14 -2242 -10
rect -2229 -14 -2206 -10
rect -2360 -34 -2356 -14
rect -2331 -18 -2328 -14
rect -2245 -18 -2242 -14
rect -2349 -22 -2328 -18
rect -2316 -22 -2260 -18
rect -2245 -22 -2221 -18
rect -2360 -38 -2345 -34
rect -2360 -58 -2356 -38
rect -2349 -46 -2328 -42
rect -2331 -50 -2312 -46
rect -2360 -62 -2345 -58
rect -2360 -82 -2356 -62
rect -2331 -66 -2328 -50
rect -2294 -54 -2290 -22
rect -2216 -34 -2206 -14
rect -2229 -38 -2206 -34
rect -2245 -46 -2221 -42
rect -2268 -50 -2242 -46
rect -2316 -58 -2260 -54
rect -2349 -70 -2328 -66
rect -2328 -79 -2304 -75
rect -2360 -86 -2345 -82
rect -2360 -106 -2356 -86
rect -2349 -94 -2328 -90
rect -2331 -106 -2328 -94
rect -2360 -110 -2345 -106
rect -2331 -110 -2312 -106
rect -2360 -130 -2356 -110
rect -2331 -114 -2328 -110
rect -2349 -118 -2328 -114
rect -2360 -134 -2345 -130
rect -2360 -154 -2356 -134
rect -2331 -138 -2328 -118
rect -2349 -142 -2328 -138
rect -2360 -158 -2345 -154
rect -2340 -158 -2328 -154
rect -2323 -158 -2312 -154
rect -2360 -182 -2356 -158
rect -2340 -162 -2337 -158
rect -2323 -162 -2320 -158
rect -2308 -159 -2304 -79
rect -2294 -111 -2290 -58
rect -2245 -66 -2242 -50
rect -2216 -58 -2206 -38
rect -2229 -62 -2206 -58
rect -2245 -70 -2221 -66
rect -2216 -82 -2206 -62
rect -2229 -86 -2206 -82
rect -2245 -94 -2221 -90
rect -2245 -106 -2242 -94
rect -2216 -106 -2206 -86
rect -2268 -110 -2242 -106
rect -2229 -110 -2206 -106
rect -2245 -114 -2242 -110
rect -2245 -118 -2221 -114
rect -2245 -138 -2242 -118
rect -2216 -130 -2206 -110
rect -2229 -134 -2206 -130
rect -2245 -142 -2221 -138
rect -2216 -154 -2206 -134
rect -2268 -158 -2253 -154
rect -2249 -158 -2233 -154
rect -2229 -158 -2206 -154
rect -2349 -166 -2337 -162
rect -2332 -166 -2320 -162
rect -2256 -162 -2253 -158
rect -2236 -162 -2233 -158
rect -2256 -166 -2241 -162
rect -2236 -166 -2221 -162
rect -2216 -182 -2206 -158
rect -2360 -186 -2252 -182
rect -2229 -186 -2206 -182
rect -2360 -197 -2356 -186
rect -2216 -197 -2206 -186
rect -2360 -201 -2345 -197
rect -2324 -201 -2206 -197
rect -2130 -595 -2126 -8
rect -2072 -8 -2057 -4
rect -2072 -28 -2068 -8
rect -2061 -16 -2040 -12
rect -2043 -28 -2040 -16
rect -2072 -32 -2057 -28
rect -2043 -32 -2024 -28
rect -2072 -52 -2068 -32
rect -2043 -36 -2040 -32
rect -2061 -40 -2040 -36
rect -2072 -56 -2057 -52
rect -2072 -76 -2068 -56
rect -2043 -60 -2040 -40
rect -2061 -64 -2040 -60
rect -2072 -80 -2057 -76
rect -2052 -80 -2040 -76
rect -2035 -80 -2024 -76
rect -2072 -104 -2068 -80
rect -2052 -84 -2049 -80
rect -2035 -84 -2032 -80
rect -2020 -81 -2016 -1
rect -2006 -33 -2002 20
rect -1957 12 -1954 28
rect -1928 20 -1918 40
rect -1941 16 -1918 20
rect -1957 8 -1933 12
rect -1928 -4 -1918 16
rect -1941 -8 -1918 -4
rect -1957 -16 -1933 -12
rect -1957 -28 -1954 -16
rect -1928 -28 -1918 -8
rect -1980 -32 -1954 -28
rect -1941 -32 -1918 -28
rect -1957 -36 -1954 -32
rect -1957 -40 -1933 -36
rect -1957 -60 -1954 -40
rect -1928 -52 -1918 -32
rect -1941 -56 -1918 -52
rect -1957 -64 -1933 -60
rect -1928 -76 -1918 -56
rect -1980 -80 -1965 -76
rect -1961 -80 -1945 -76
rect -1941 -80 -1918 -76
rect -2061 -88 -2049 -84
rect -2044 -88 -2032 -84
rect -1968 -84 -1965 -80
rect -1948 -84 -1945 -80
rect -1968 -88 -1953 -84
rect -1948 -88 -1933 -84
rect -1928 -104 -1918 -80
rect -2072 -108 -1964 -104
rect -1941 -108 -1918 -104
rect -2072 -119 -2068 -108
rect -1928 -119 -1918 -108
rect -2103 -123 -2057 -119
rect -2036 -123 -1918 -119
rect -1848 148 -1765 152
rect -2103 -352 -2099 -123
rect -1953 -346 -1949 -123
rect -1959 -352 -1949 -346
rect -2103 -356 -2088 -352
rect -2074 -356 -2055 -352
rect -2011 -356 -1985 -352
rect -1972 -356 -1949 -352
rect -2103 -376 -2099 -356
rect -2074 -360 -2071 -356
rect -1988 -360 -1985 -356
rect -2092 -364 -2071 -360
rect -2059 -364 -2003 -360
rect -1988 -364 -1964 -360
rect -2103 -380 -2088 -376
rect -2103 -400 -2099 -380
rect -2092 -388 -2071 -384
rect -2074 -392 -2055 -388
rect -2103 -404 -2088 -400
rect -2103 -424 -2099 -404
rect -2074 -408 -2071 -392
rect -2037 -396 -2033 -364
rect -1959 -376 -1949 -356
rect -1972 -380 -1949 -376
rect -1988 -388 -1964 -384
rect -2011 -392 -1985 -388
rect -2059 -400 -2003 -396
rect -2092 -412 -2071 -408
rect -2071 -421 -2047 -417
rect -2103 -428 -2088 -424
rect -2103 -448 -2099 -428
rect -2092 -436 -2071 -432
rect -2074 -448 -2071 -436
rect -2103 -452 -2088 -448
rect -2074 -452 -2055 -448
rect -2103 -472 -2099 -452
rect -2074 -456 -2071 -452
rect -2092 -460 -2071 -456
rect -2103 -476 -2088 -472
rect -2103 -496 -2099 -476
rect -2074 -480 -2071 -460
rect -2092 -484 -2071 -480
rect -2103 -500 -2088 -496
rect -2083 -500 -2071 -496
rect -2066 -500 -2055 -496
rect -2103 -524 -2099 -500
rect -2083 -504 -2080 -500
rect -2066 -504 -2063 -500
rect -2051 -501 -2047 -421
rect -2037 -453 -2033 -400
rect -1988 -408 -1985 -392
rect -1959 -400 -1949 -380
rect -1972 -404 -1949 -400
rect -1988 -412 -1964 -408
rect -1959 -424 -1949 -404
rect -1848 -413 -1844 148
rect -1824 133 -1677 137
rect -1834 109 -1781 113
rect -1798 94 -1644 98
rect -1720 69 -1658 73
rect -1720 48 -1716 69
rect -1674 48 -1670 54
rect -1720 44 -1708 48
rect -1690 44 -1670 48
rect -1747 21 -1741 32
rect -1763 17 -1741 21
rect -1810 5 -1802 9
rect -1814 -20 -1810 5
rect -1747 -1 -1741 17
rect -1763 -5 -1741 -1
rect -1747 -20 -1741 -5
rect -1814 -24 -1784 -20
rect -1763 -24 -1741 -20
rect -1814 -43 -1810 -24
rect -1747 -33 -1741 -24
rect -1720 3 -1716 44
rect -1712 36 -1682 40
rect -1703 24 -1699 36
rect -1703 20 -1688 24
rect -1720 -1 -1705 3
rect -1720 -24 -1716 -1
rect -1720 -28 -1705 -24
rect -1720 -43 -1716 -28
rect -1814 -48 -1716 -43
rect -1692 -47 -1688 20
rect -1814 -59 -1810 -48
rect -1829 -63 -1810 -59
rect -1829 -172 -1825 -63
rect -1674 -78 -1670 44
rect -1662 47 -1658 69
rect -1615 47 -1611 159
rect -1362 135 -1358 150
rect -1398 131 -1358 135
rect -1662 43 -1649 47
rect -1631 43 -1611 47
rect -1662 31 -1658 43
rect -1653 35 -1623 39
rect -1644 -26 -1640 35
rect -1615 4 -1611 43
rect -1632 0 -1611 4
rect -1615 -30 -1611 0
rect -1632 -34 -1611 -30
rect -1741 -79 -1670 -78
rect -1615 -79 -1611 -34
rect -1741 -83 -1611 -79
rect -1419 -77 -1414 127
rect -1398 84 -1394 131
rect -1382 84 -1228 88
rect -1304 59 -1242 63
rect -1304 38 -1300 59
rect -1258 38 -1254 44
rect -1304 34 -1292 38
rect -1274 34 -1254 38
rect -1331 11 -1325 22
rect -1347 7 -1325 11
rect -1394 -5 -1386 -1
rect -1398 -30 -1394 -5
rect -1331 -11 -1325 7
rect -1347 -15 -1325 -11
rect -1331 -30 -1325 -15
rect -1398 -34 -1368 -30
rect -1347 -34 -1325 -30
rect -1398 -53 -1394 -34
rect -1331 -43 -1325 -34
rect -1304 -7 -1300 34
rect -1296 26 -1266 30
rect -1287 14 -1283 26
rect -1287 10 -1272 14
rect -1304 -11 -1289 -7
rect -1304 -34 -1300 -11
rect -1304 -38 -1289 -34
rect -1304 -53 -1300 -38
rect -1398 -58 -1300 -53
rect -1276 -57 -1272 10
rect -1616 -166 -1611 -83
rect -1398 -85 -1394 -58
rect -1685 -170 -1611 -166
rect -1578 -89 -1394 -85
rect -1258 -88 -1254 34
rect -1246 37 -1242 59
rect -1199 37 -1195 159
rect -934 117 -780 121
rect -1137 100 -1066 104
rect -856 92 -794 96
rect -856 71 -852 92
rect -810 71 -806 77
rect -856 67 -844 71
rect -826 67 -806 71
rect -883 44 -877 55
rect -899 40 -877 44
rect -1246 33 -1233 37
rect -1215 33 -1195 37
rect -1246 21 -1242 33
rect -1237 25 -1207 29
rect -1228 -36 -1224 25
rect -1199 -6 -1195 33
rect -1216 -10 -1195 -6
rect -1199 -40 -1195 -10
rect -946 28 -938 32
rect -950 3 -946 28
rect -883 22 -877 40
rect -899 18 -877 22
rect -883 3 -877 18
rect -950 -1 -920 3
rect -899 -1 -877 3
rect -950 -20 -946 -1
rect -883 -10 -877 -1
rect -856 26 -852 67
rect -848 59 -818 63
rect -839 47 -835 59
rect -839 43 -824 47
rect -856 22 -841 26
rect -856 -1 -852 22
rect -856 -5 -841 -1
rect -856 -20 -852 -5
rect -950 -25 -852 -20
rect -828 -24 -824 43
rect -950 -36 -946 -25
rect -1216 -44 -1195 -40
rect -1578 -132 -1574 -89
rect -1325 -89 -1254 -88
rect -1199 -89 -1195 -44
rect -1325 -93 -1195 -89
rect -1419 -114 -1414 -98
rect -1199 -126 -1195 -93
rect -1434 -130 -1195 -126
rect -1160 -40 -946 -36
rect -1160 -83 -1156 -40
rect -810 -55 -806 67
rect -798 70 -794 92
rect -751 70 -747 159
rect -798 66 -785 70
rect -767 66 -747 70
rect -798 54 -794 66
rect -789 58 -759 62
rect -780 -3 -776 58
rect -751 27 -747 66
rect -768 23 -747 27
rect -751 -7 -747 23
rect -768 -11 -747 -7
rect -877 -56 -806 -55
rect -751 -56 -747 -11
rect -877 -60 -747 -56
rect -752 -77 -747 -60
rect -1016 -81 -747 -77
rect -1016 -83 -1006 -81
rect -1160 -87 -1145 -83
rect -1131 -87 -1112 -83
rect -1068 -87 -1042 -83
rect -1029 -87 -1006 -83
rect -1160 -107 -1156 -87
rect -1131 -91 -1128 -87
rect -1045 -91 -1042 -87
rect -1149 -95 -1128 -91
rect -1116 -95 -1060 -91
rect -1045 -95 -1021 -91
rect -1160 -111 -1145 -107
rect -1434 -132 -1424 -130
rect -1578 -136 -1563 -132
rect -1549 -136 -1530 -132
rect -1486 -136 -1460 -132
rect -1447 -136 -1424 -132
rect -1578 -156 -1574 -136
rect -1549 -140 -1546 -136
rect -1463 -140 -1460 -136
rect -1567 -144 -1546 -140
rect -1534 -144 -1478 -140
rect -1463 -144 -1439 -140
rect -1578 -160 -1563 -156
rect -1685 -172 -1675 -170
rect -1829 -176 -1814 -172
rect -1800 -176 -1781 -172
rect -1737 -176 -1711 -172
rect -1698 -176 -1675 -172
rect -1829 -196 -1825 -176
rect -1800 -180 -1797 -176
rect -1714 -180 -1711 -176
rect -1818 -184 -1797 -180
rect -1785 -184 -1729 -180
rect -1714 -184 -1690 -180
rect -1829 -200 -1814 -196
rect -1829 -220 -1825 -200
rect -1818 -208 -1797 -204
rect -1800 -212 -1781 -208
rect -1829 -224 -1814 -220
rect -1829 -244 -1825 -224
rect -1800 -228 -1797 -212
rect -1763 -216 -1759 -184
rect -1685 -196 -1675 -176
rect -1698 -200 -1675 -196
rect -1714 -208 -1690 -204
rect -1737 -212 -1711 -208
rect -1785 -220 -1729 -216
rect -1818 -232 -1797 -228
rect -1797 -241 -1773 -237
rect -1829 -248 -1814 -244
rect -1829 -268 -1825 -248
rect -1818 -256 -1797 -252
rect -1800 -268 -1797 -256
rect -1829 -272 -1814 -268
rect -1800 -272 -1781 -268
rect -1829 -292 -1825 -272
rect -1800 -276 -1797 -272
rect -1818 -280 -1797 -276
rect -1829 -296 -1814 -292
rect -1829 -316 -1825 -296
rect -1800 -300 -1797 -280
rect -1818 -304 -1797 -300
rect -1829 -320 -1814 -316
rect -1809 -320 -1797 -316
rect -1792 -320 -1781 -316
rect -1829 -344 -1825 -320
rect -1809 -324 -1806 -320
rect -1792 -324 -1789 -320
rect -1777 -321 -1773 -241
rect -1763 -273 -1759 -220
rect -1714 -228 -1711 -212
rect -1685 -220 -1675 -200
rect -1698 -224 -1675 -220
rect -1714 -232 -1690 -228
rect -1685 -244 -1675 -224
rect -1698 -248 -1675 -244
rect -1714 -256 -1690 -252
rect -1714 -268 -1711 -256
rect -1685 -268 -1675 -248
rect -1737 -272 -1711 -268
rect -1698 -272 -1675 -268
rect -1714 -276 -1711 -272
rect -1714 -280 -1690 -276
rect -1714 -300 -1711 -280
rect -1685 -292 -1675 -272
rect -1698 -296 -1675 -292
rect -1714 -304 -1690 -300
rect -1685 -316 -1675 -296
rect -1737 -320 -1722 -316
rect -1718 -320 -1702 -316
rect -1698 -320 -1675 -316
rect -1818 -328 -1806 -324
rect -1801 -328 -1789 -324
rect -1725 -324 -1722 -320
rect -1705 -324 -1702 -320
rect -1725 -328 -1710 -324
rect -1705 -328 -1690 -324
rect -1685 -344 -1675 -320
rect -1578 -180 -1574 -160
rect -1567 -168 -1546 -164
rect -1549 -172 -1530 -168
rect -1578 -184 -1563 -180
rect -1578 -204 -1574 -184
rect -1549 -188 -1546 -172
rect -1512 -176 -1508 -144
rect -1434 -156 -1424 -136
rect -1447 -160 -1424 -156
rect -1463 -168 -1439 -164
rect -1486 -172 -1460 -168
rect -1534 -180 -1478 -176
rect -1567 -192 -1546 -188
rect -1546 -201 -1522 -197
rect -1578 -208 -1563 -204
rect -1578 -228 -1574 -208
rect -1567 -216 -1546 -212
rect -1549 -228 -1546 -216
rect -1578 -232 -1563 -228
rect -1549 -232 -1530 -228
rect -1578 -252 -1574 -232
rect -1549 -236 -1546 -232
rect -1567 -240 -1546 -236
rect -1578 -256 -1563 -252
rect -1578 -276 -1574 -256
rect -1549 -260 -1546 -240
rect -1567 -264 -1546 -260
rect -1578 -280 -1563 -276
rect -1558 -280 -1546 -276
rect -1541 -280 -1530 -276
rect -1578 -304 -1574 -280
rect -1558 -284 -1555 -280
rect -1541 -284 -1538 -280
rect -1526 -281 -1522 -201
rect -1512 -233 -1508 -180
rect -1463 -188 -1460 -172
rect -1434 -180 -1424 -160
rect -1447 -184 -1424 -180
rect -1463 -192 -1439 -188
rect -1434 -204 -1424 -184
rect -1447 -208 -1424 -204
rect -1463 -216 -1439 -212
rect -1463 -228 -1460 -216
rect -1434 -228 -1424 -208
rect -1486 -232 -1460 -228
rect -1447 -232 -1424 -228
rect -1463 -236 -1460 -232
rect -1463 -240 -1439 -236
rect -1463 -260 -1460 -240
rect -1434 -252 -1424 -232
rect -1447 -256 -1424 -252
rect -1463 -264 -1439 -260
rect -1434 -276 -1424 -256
rect -1160 -131 -1156 -111
rect -1149 -119 -1128 -115
rect -1131 -123 -1112 -119
rect -1160 -135 -1145 -131
rect -1160 -155 -1156 -135
rect -1131 -139 -1128 -123
rect -1094 -127 -1090 -95
rect -1016 -107 -1006 -87
rect -1029 -111 -1006 -107
rect -1045 -119 -1021 -115
rect -1068 -123 -1042 -119
rect -1116 -131 -1060 -127
rect -1149 -143 -1128 -139
rect -1128 -152 -1104 -148
rect -1160 -159 -1145 -155
rect -1160 -179 -1156 -159
rect -1149 -167 -1128 -163
rect -1131 -179 -1128 -167
rect -1160 -183 -1145 -179
rect -1131 -183 -1112 -179
rect -1160 -203 -1156 -183
rect -1131 -187 -1128 -183
rect -1149 -191 -1128 -187
rect -1160 -207 -1145 -203
rect -1160 -227 -1156 -207
rect -1131 -211 -1128 -191
rect -1149 -215 -1128 -211
rect -1160 -231 -1145 -227
rect -1140 -231 -1128 -227
rect -1123 -231 -1112 -227
rect -1160 -255 -1156 -231
rect -1140 -235 -1137 -231
rect -1123 -235 -1120 -231
rect -1108 -232 -1104 -152
rect -1094 -184 -1090 -131
rect -1045 -139 -1042 -123
rect -1016 -131 -1006 -111
rect -1029 -135 -1006 -131
rect -1045 -143 -1021 -139
rect -1016 -155 -1006 -135
rect -1029 -159 -1006 -155
rect -1045 -167 -1021 -163
rect -1045 -179 -1042 -167
rect -1016 -179 -1006 -159
rect -1068 -183 -1042 -179
rect -1029 -183 -1006 -179
rect -1045 -187 -1042 -183
rect -1045 -191 -1021 -187
rect -1045 -211 -1042 -191
rect -1016 -203 -1006 -183
rect -1029 -207 -1006 -203
rect -1045 -215 -1021 -211
rect -1016 -227 -1006 -207
rect -1068 -231 -1053 -227
rect -1049 -231 -1033 -227
rect -1029 -231 -1006 -227
rect -1149 -239 -1137 -235
rect -1132 -239 -1120 -235
rect -1056 -235 -1053 -231
rect -1036 -235 -1033 -231
rect -1056 -239 -1041 -235
rect -1036 -239 -1021 -235
rect -1016 -255 -1006 -231
rect -1160 -259 -1052 -255
rect -1029 -259 -1006 -255
rect -1160 -270 -1156 -259
rect -1016 -270 -1006 -259
rect -1160 -272 -1145 -270
rect -1486 -280 -1471 -276
rect -1467 -280 -1451 -276
rect -1447 -280 -1424 -276
rect -1567 -288 -1555 -284
rect -1550 -288 -1538 -284
rect -1474 -284 -1471 -280
rect -1454 -284 -1451 -280
rect -1474 -288 -1459 -284
rect -1454 -288 -1439 -284
rect -1434 -304 -1424 -280
rect -1578 -308 -1470 -304
rect -1447 -308 -1424 -304
rect -1578 -319 -1574 -308
rect -1434 -319 -1424 -308
rect -1574 -323 -1563 -319
rect -1542 -323 -1424 -319
rect -1377 -274 -1145 -272
rect -1124 -274 -1006 -270
rect -1377 -276 -1156 -274
rect -1377 -319 -1373 -276
rect -1082 -313 -1078 -274
rect -1233 -317 -1078 -313
rect -1233 -319 -1223 -317
rect -1377 -323 -1362 -319
rect -1348 -323 -1329 -319
rect -1285 -323 -1259 -319
rect -1246 -323 -1223 -319
rect -1829 -348 -1721 -344
rect -1698 -348 -1675 -344
rect -1829 -359 -1825 -348
rect -1685 -359 -1675 -348
rect -1836 -363 -1814 -359
rect -1793 -363 -1675 -359
rect -1664 -355 -1557 -351
rect -1972 -428 -1949 -424
rect -1988 -436 -1964 -432
rect -1988 -448 -1985 -436
rect -1959 -448 -1949 -428
rect -2011 -452 -1985 -448
rect -1972 -452 -1949 -448
rect -1988 -456 -1985 -452
rect -1988 -460 -1964 -456
rect -1988 -480 -1985 -460
rect -1959 -472 -1949 -452
rect -1972 -476 -1949 -472
rect -1988 -484 -1964 -480
rect -1959 -496 -1949 -476
rect -2011 -500 -1996 -496
rect -1992 -500 -1976 -496
rect -1972 -500 -1949 -496
rect -2092 -508 -2080 -504
rect -2075 -508 -2063 -504
rect -1999 -504 -1996 -500
rect -1979 -504 -1976 -500
rect -1999 -508 -1984 -504
rect -1979 -508 -1964 -504
rect -1959 -524 -1949 -500
rect -2103 -528 -1995 -524
rect -1972 -528 -1949 -524
rect -2103 -539 -2099 -528
rect -1959 -539 -1949 -528
rect -2103 -543 -2088 -539
rect -2067 -543 -1949 -539
rect -1836 -472 -1832 -363
rect -1686 -466 -1682 -363
rect -1664 -446 -1660 -355
rect -1648 -388 -1531 -384
rect -1648 -456 -1644 -388
rect -1535 -390 -1531 -388
rect -1630 -403 -1476 -399
rect -1692 -472 -1682 -466
rect -1836 -476 -1821 -472
rect -1807 -476 -1788 -472
rect -1744 -476 -1718 -472
rect -1705 -476 -1682 -472
rect -1836 -496 -1832 -476
rect -1807 -480 -1804 -476
rect -1721 -480 -1718 -476
rect -1825 -484 -1804 -480
rect -1792 -484 -1736 -480
rect -1721 -484 -1697 -480
rect -1836 -500 -1821 -496
rect -1836 -520 -1832 -500
rect -1825 -508 -1804 -504
rect -1807 -512 -1788 -508
rect -1836 -524 -1821 -520
rect -1956 -595 -1952 -543
rect -2130 -599 -1952 -595
rect -1836 -544 -1832 -524
rect -1807 -528 -1804 -512
rect -1770 -516 -1766 -484
rect -1692 -496 -1682 -476
rect -1705 -500 -1682 -496
rect -1721 -508 -1697 -504
rect -1744 -512 -1718 -508
rect -1792 -520 -1736 -516
rect -1825 -532 -1804 -528
rect -1804 -541 -1780 -537
rect -1836 -548 -1821 -544
rect -1836 -568 -1832 -548
rect -1825 -556 -1804 -552
rect -1807 -568 -1804 -556
rect -1836 -572 -1821 -568
rect -1807 -572 -1788 -568
rect -1836 -592 -1832 -572
rect -1807 -576 -1804 -572
rect -1825 -580 -1804 -576
rect -1836 -596 -1821 -592
rect -1836 -616 -1832 -596
rect -1807 -600 -1804 -580
rect -1825 -604 -1804 -600
rect -1836 -620 -1821 -616
rect -1816 -620 -1804 -616
rect -1799 -620 -1788 -616
rect -1836 -644 -1832 -620
rect -1816 -624 -1813 -620
rect -1799 -624 -1796 -620
rect -1784 -621 -1780 -541
rect -1770 -573 -1766 -520
rect -1721 -528 -1718 -512
rect -1692 -520 -1682 -500
rect -1705 -524 -1682 -520
rect -1721 -532 -1697 -528
rect -1692 -544 -1682 -524
rect -1705 -548 -1682 -544
rect -1721 -556 -1697 -552
rect -1721 -568 -1718 -556
rect -1692 -568 -1682 -548
rect -1744 -572 -1718 -568
rect -1705 -572 -1682 -568
rect -1721 -576 -1718 -572
rect -1721 -580 -1697 -576
rect -1721 -600 -1718 -580
rect -1692 -592 -1682 -572
rect -1705 -596 -1682 -592
rect -1721 -604 -1697 -600
rect -1692 -616 -1682 -596
rect -1744 -620 -1729 -616
rect -1725 -620 -1709 -616
rect -1705 -620 -1682 -616
rect -1825 -628 -1813 -624
rect -1808 -628 -1796 -624
rect -1732 -624 -1729 -620
rect -1712 -624 -1709 -620
rect -1732 -628 -1717 -624
rect -1712 -628 -1697 -624
rect -1692 -644 -1682 -620
rect -1836 -648 -1728 -644
rect -1705 -648 -1682 -644
rect -1836 -659 -1832 -648
rect -1692 -659 -1682 -648
rect -1836 -663 -1821 -659
rect -1800 -663 -1682 -659
rect -1660 -460 -1644 -456
rect -1552 -428 -1490 -424
rect -1552 -449 -1548 -428
rect -1506 -449 -1502 -443
rect -1552 -453 -1540 -449
rect -1522 -453 -1502 -449
rect -1660 -684 -1656 -460
rect -1579 -476 -1573 -465
rect -1595 -480 -1573 -476
rect -1642 -492 -1634 -488
rect -1646 -517 -1642 -492
rect -1579 -498 -1573 -480
rect -1595 -502 -1573 -498
rect -1579 -517 -1573 -502
rect -1646 -521 -1616 -517
rect -1595 -521 -1573 -517
rect -1646 -540 -1642 -521
rect -1579 -530 -1573 -521
rect -1552 -494 -1548 -453
rect -1544 -461 -1514 -457
rect -1535 -473 -1531 -461
rect -1535 -477 -1520 -473
rect -1552 -498 -1537 -494
rect -1552 -521 -1548 -498
rect -1552 -525 -1537 -521
rect -1552 -540 -1548 -525
rect -1646 -545 -1548 -540
rect -1524 -544 -1520 -477
rect -1506 -575 -1502 -453
rect -1494 -450 -1490 -428
rect -1447 -450 -1443 -323
rect -1494 -454 -1481 -450
rect -1463 -454 -1443 -450
rect -1494 -466 -1490 -454
rect -1485 -462 -1455 -458
rect -1476 -523 -1472 -462
rect -1447 -493 -1443 -454
rect -1464 -497 -1443 -493
rect -1447 -527 -1443 -497
rect -1377 -343 -1373 -323
rect -1348 -327 -1345 -323
rect -1262 -327 -1259 -323
rect -1366 -331 -1345 -327
rect -1333 -331 -1277 -327
rect -1262 -331 -1238 -327
rect -1377 -347 -1362 -343
rect -1377 -367 -1373 -347
rect -1366 -355 -1345 -351
rect -1348 -359 -1329 -355
rect -1377 -371 -1362 -367
rect -1377 -391 -1373 -371
rect -1348 -375 -1345 -359
rect -1311 -363 -1307 -331
rect -1233 -343 -1223 -323
rect -1246 -347 -1223 -343
rect -1262 -355 -1238 -351
rect -1285 -359 -1259 -355
rect -1333 -367 -1277 -363
rect -1366 -379 -1345 -375
rect -1345 -388 -1321 -384
rect -1377 -395 -1362 -391
rect -1377 -415 -1373 -395
rect -1366 -403 -1345 -399
rect -1348 -415 -1345 -403
rect -1377 -419 -1362 -415
rect -1348 -419 -1329 -415
rect -1377 -439 -1373 -419
rect -1348 -423 -1345 -419
rect -1366 -427 -1345 -423
rect -1377 -443 -1362 -439
rect -1377 -463 -1373 -443
rect -1348 -447 -1345 -427
rect -1366 -451 -1345 -447
rect -1377 -467 -1362 -463
rect -1357 -467 -1345 -463
rect -1340 -467 -1329 -463
rect -1377 -491 -1373 -467
rect -1357 -471 -1354 -467
rect -1340 -471 -1337 -467
rect -1325 -468 -1321 -388
rect -1311 -420 -1307 -367
rect -1262 -375 -1259 -359
rect -1233 -367 -1223 -347
rect -1246 -371 -1223 -367
rect -1262 -379 -1238 -375
rect -1233 -391 -1223 -371
rect -1246 -395 -1223 -391
rect -1262 -403 -1238 -399
rect -1262 -415 -1259 -403
rect -1233 -415 -1223 -395
rect -1285 -419 -1259 -415
rect -1246 -419 -1223 -415
rect -1262 -423 -1259 -419
rect -1262 -427 -1238 -423
rect -1262 -447 -1259 -427
rect -1233 -439 -1223 -419
rect -1246 -443 -1223 -439
rect -1262 -451 -1238 -447
rect -1233 -463 -1223 -443
rect -1285 -467 -1270 -463
rect -1266 -467 -1250 -463
rect -1246 -467 -1223 -463
rect -1366 -475 -1354 -471
rect -1349 -475 -1337 -471
rect -1273 -471 -1270 -467
rect -1253 -471 -1250 -467
rect -1273 -475 -1258 -471
rect -1253 -475 -1238 -471
rect -1233 -491 -1223 -467
rect -1377 -495 -1269 -491
rect -1246 -495 -1223 -491
rect -1377 -506 -1373 -495
rect -1233 -506 -1223 -495
rect -1377 -510 -1362 -506
rect -1341 -510 -1223 -506
rect -1464 -531 -1443 -527
rect -1573 -576 -1502 -575
rect -1447 -576 -1443 -531
rect -1573 -580 -1443 -576
rect -1717 -688 -1656 -684
<< ntransistor >>
rect -2060 207 -2056 209
rect -2043 207 -2039 209
rect -1971 206 -1967 208
rect -1954 206 -1950 208
rect -1884 206 -1880 208
rect -1867 206 -1863 208
rect -1795 207 -1791 209
rect -1778 207 -1774 209
rect -1707 207 -1703 209
rect -1690 207 -1686 209
rect -1617 207 -1613 209
rect -1600 207 -1596 209
rect -1525 207 -1521 209
rect -1508 207 -1504 209
rect -1430 207 -1426 209
rect -1413 207 -1409 209
rect -1341 207 -1337 209
rect -1324 207 -1320 209
rect -1249 208 -1245 210
rect -1232 208 -1228 210
rect -1155 207 -1151 209
rect -1138 207 -1134 209
rect -1067 207 -1063 209
rect -1050 207 -1046 209
rect -977 207 -973 209
rect -960 207 -956 209
rect -886 207 -882 209
rect -869 207 -865 209
rect -795 207 -791 209
rect -778 207 -774 209
rect -706 207 -702 209
rect -689 207 -685 209
rect -2042 178 -2038 180
rect -1953 177 -1949 179
rect -1866 177 -1862 179
rect -1777 178 -1773 180
rect -1689 178 -1685 180
rect -1599 178 -1595 180
rect -1507 178 -1503 180
rect -1412 178 -1408 180
rect -1323 178 -1319 180
rect -1231 179 -1227 181
rect -1137 178 -1133 180
rect -1049 178 -1045 180
rect -959 178 -955 180
rect -868 178 -864 180
rect -777 178 -773 180
rect -688 178 -684 180
rect -848 64 -844 66
rect -2061 61 -2057 63
rect -2028 61 -2024 63
rect -789 63 -785 65
rect -1712 41 -1708 43
rect -2061 37 -2057 39
rect -1653 40 -1649 42
rect -1296 31 -1292 33
rect -2028 25 -2024 27
rect -1237 30 -1233 32
rect -2061 13 -2057 15
rect -2061 -11 -2057 -9
rect -2349 -17 -2345 -15
rect -2316 -17 -2312 -15
rect -1806 2 -1802 4
rect -1789 2 -1785 4
rect -942 25 -938 27
rect -925 25 -921 27
rect -845 19 -841 21
rect -823 20 -819 22
rect -1709 -4 -1705 -2
rect -1687 -3 -1683 -1
rect -1788 -27 -1784 -25
rect -2061 -35 -2057 -33
rect -2028 -35 -2024 -33
rect -2349 -41 -2345 -39
rect -2316 -53 -2312 -51
rect -2061 -59 -2057 -57
rect -2349 -65 -2345 -63
rect -1390 -8 -1386 -6
rect -1373 -8 -1369 -6
rect -924 -4 -920 -2
rect -1293 -14 -1289 -12
rect -1271 -13 -1267 -11
rect -1709 -31 -1705 -29
rect -1687 -30 -1683 -28
rect -1372 -37 -1368 -35
rect -1293 -41 -1289 -39
rect -1271 -40 -1267 -38
rect -845 -8 -841 -6
rect -823 -7 -819 -5
rect -2061 -83 -2057 -81
rect -2044 -83 -2040 -81
rect -2028 -83 -2024 -81
rect -2349 -89 -2345 -87
rect -1149 -90 -1145 -88
rect -1116 -90 -1112 -88
rect -1968 -111 -1964 -109
rect -2349 -113 -2345 -111
rect -2316 -113 -2312 -111
rect -1149 -114 -1145 -112
rect -2061 -126 -2057 -124
rect -1116 -126 -1112 -124
rect -2349 -137 -2345 -135
rect -1567 -139 -1563 -137
rect -1534 -139 -1530 -137
rect -1149 -138 -1145 -136
rect -2349 -161 -2345 -159
rect -2332 -161 -2328 -159
rect -2316 -161 -2312 -159
rect -1567 -163 -1563 -161
rect -1149 -162 -1145 -160
rect -1534 -175 -1530 -173
rect -1818 -179 -1814 -177
rect -1785 -179 -1781 -177
rect -1567 -187 -1563 -185
rect -1149 -186 -1145 -184
rect -1116 -186 -1112 -184
rect -2256 -189 -2252 -187
rect -2349 -204 -2345 -202
rect -1818 -203 -1814 -201
rect -1567 -211 -1563 -209
rect -1149 -210 -1145 -208
rect -1785 -215 -1781 -213
rect -1818 -227 -1814 -225
rect -1567 -235 -1563 -233
rect -1534 -235 -1530 -233
rect -1149 -234 -1145 -232
rect -1132 -234 -1128 -232
rect -1116 -234 -1112 -232
rect -1818 -251 -1814 -249
rect -1567 -259 -1563 -257
rect -1056 -262 -1052 -260
rect -1818 -275 -1814 -273
rect -1785 -275 -1781 -273
rect -1149 -277 -1145 -275
rect -1567 -283 -1563 -281
rect -1550 -283 -1546 -281
rect -1534 -283 -1530 -281
rect -1818 -299 -1814 -297
rect -1474 -311 -1470 -309
rect -1818 -323 -1814 -321
rect -1801 -323 -1797 -321
rect -1785 -323 -1781 -321
rect -1567 -326 -1563 -324
rect -1366 -326 -1362 -324
rect -1333 -326 -1329 -324
rect -1725 -351 -1721 -349
rect -1366 -350 -1362 -348
rect -2092 -359 -2088 -357
rect -2059 -359 -2055 -357
rect -1333 -362 -1329 -360
rect -1818 -366 -1814 -364
rect -1366 -374 -1362 -372
rect -2092 -383 -2088 -381
rect -2059 -395 -2055 -393
rect -1366 -398 -1362 -396
rect -2092 -407 -2088 -405
rect -1366 -422 -1362 -420
rect -1333 -422 -1329 -420
rect -2092 -431 -2088 -429
rect -1366 -446 -1362 -444
rect -2092 -455 -2088 -453
rect -2059 -455 -2055 -453
rect -1544 -456 -1540 -454
rect -1485 -457 -1481 -455
rect -1366 -470 -1362 -468
rect -1349 -470 -1345 -468
rect -1333 -470 -1329 -468
rect -2092 -479 -2088 -477
rect -1825 -479 -1821 -477
rect -1792 -479 -1788 -477
rect -2092 -503 -2088 -501
rect -2075 -503 -2071 -501
rect -2059 -503 -2055 -501
rect -1825 -503 -1821 -501
rect -1638 -495 -1634 -493
rect -1621 -495 -1617 -493
rect -1273 -498 -1269 -496
rect -1541 -501 -1537 -499
rect -1519 -500 -1515 -498
rect -1792 -515 -1788 -513
rect -1620 -524 -1616 -522
rect -1825 -527 -1821 -525
rect -1999 -531 -1995 -529
rect -2092 -546 -2088 -544
rect -1825 -551 -1821 -549
rect -1366 -513 -1362 -511
rect -1541 -528 -1537 -526
rect -1519 -527 -1515 -525
rect -1825 -575 -1821 -573
rect -1792 -575 -1788 -573
rect -1825 -599 -1821 -597
rect -1825 -623 -1821 -621
rect -1808 -623 -1804 -621
rect -1792 -623 -1788 -621
rect -1732 -651 -1728 -649
rect -1825 -666 -1821 -664
<< ptransistor >>
rect -2017 219 -2009 221
rect -2017 197 -2009 199
rect -1928 218 -1920 220
rect -1928 196 -1920 198
rect -1841 218 -1833 220
rect -1841 196 -1833 198
rect -1752 219 -1744 221
rect -1752 197 -1744 199
rect -1664 219 -1656 221
rect -1664 197 -1656 199
rect -1574 219 -1566 221
rect -1574 197 -1566 199
rect -1482 219 -1474 221
rect -1482 197 -1474 199
rect -1387 219 -1379 221
rect -1387 197 -1379 199
rect -1298 219 -1290 221
rect -1298 197 -1290 199
rect -1206 220 -1198 222
rect -1206 198 -1198 200
rect -1112 219 -1104 221
rect -1112 197 -1104 199
rect -1024 219 -1016 221
rect -1024 197 -1016 199
rect -934 219 -926 221
rect -934 197 -926 199
rect -843 219 -835 221
rect -843 197 -835 199
rect -752 219 -744 221
rect -752 197 -744 199
rect -663 219 -655 221
rect -663 197 -655 199
rect -2017 178 -2009 180
rect -1928 177 -1920 179
rect -1841 177 -1833 179
rect -1752 178 -1744 180
rect -1664 178 -1656 180
rect -1574 178 -1566 180
rect -1482 178 -1474 180
rect -1387 178 -1379 180
rect -1298 178 -1290 180
rect -1206 179 -1199 181
rect -1112 178 -1104 180
rect -1024 178 -1016 180
rect -934 178 -926 180
rect -843 178 -835 180
rect -752 178 -744 180
rect -663 178 -655 180
rect -826 64 -818 66
rect -1980 61 -1972 63
rect -1941 61 -1933 63
rect -767 63 -759 65
rect -1690 41 -1682 43
rect -1941 37 -1933 39
rect -1631 40 -1623 42
rect -1274 31 -1266 33
rect -1980 25 -1972 27
rect -1215 30 -1207 32
rect -1941 13 -1933 15
rect -1941 -11 -1933 -9
rect -2268 -17 -2260 -15
rect -2229 -17 -2221 -15
rect -1763 14 -1755 16
rect -899 37 -891 39
rect -794 20 -786 22
rect -768 20 -760 22
rect -899 15 -891 17
rect -1658 -3 -1650 -1
rect -1632 -3 -1624 -1
rect -1763 -8 -1755 -6
rect -1763 -27 -1755 -25
rect -1980 -35 -1972 -33
rect -1941 -35 -1933 -33
rect -2229 -41 -2221 -39
rect -2268 -53 -2260 -51
rect -1941 -59 -1933 -57
rect -2229 -65 -2221 -63
rect -1347 4 -1339 6
rect -899 -4 -891 -2
rect -1242 -13 -1234 -11
rect -1216 -13 -1208 -11
rect -1347 -18 -1339 -16
rect -1658 -37 -1650 -35
rect -1632 -37 -1624 -35
rect -1347 -37 -1339 -35
rect -794 -14 -786 -12
rect -768 -14 -760 -12
rect -1242 -47 -1234 -45
rect -1216 -47 -1208 -45
rect -1980 -83 -1972 -81
rect -1961 -83 -1953 -81
rect -1941 -83 -1933 -81
rect -2229 -89 -2221 -87
rect -1068 -90 -1060 -88
rect -1029 -90 -1021 -88
rect -1941 -111 -1933 -109
rect -2268 -113 -2260 -111
rect -2229 -113 -2221 -111
rect -1029 -114 -1021 -112
rect -2036 -126 -2028 -124
rect -1068 -126 -1060 -124
rect -2229 -137 -2221 -135
rect -1486 -139 -1478 -137
rect -1447 -139 -1439 -137
rect -1029 -138 -1021 -136
rect -2268 -161 -2260 -159
rect -2249 -161 -2241 -159
rect -2229 -161 -2221 -159
rect -1447 -163 -1439 -161
rect -1029 -162 -1021 -160
rect -1486 -175 -1478 -173
rect -1737 -179 -1729 -177
rect -1698 -179 -1690 -177
rect -1447 -187 -1439 -185
rect -1068 -186 -1060 -184
rect -1029 -186 -1021 -184
rect -2229 -189 -2221 -187
rect -2324 -204 -2316 -202
rect -1698 -203 -1690 -201
rect -1447 -211 -1439 -209
rect -1029 -210 -1021 -208
rect -1737 -215 -1729 -213
rect -1698 -227 -1690 -225
rect -1486 -235 -1478 -233
rect -1447 -235 -1439 -233
rect -1068 -234 -1060 -232
rect -1049 -234 -1041 -232
rect -1029 -234 -1021 -232
rect -1698 -251 -1690 -249
rect -1447 -259 -1439 -257
rect -1029 -262 -1021 -260
rect -1737 -275 -1729 -273
rect -1698 -275 -1690 -273
rect -1124 -277 -1116 -275
rect -1486 -283 -1478 -281
rect -1467 -283 -1459 -281
rect -1447 -283 -1439 -281
rect -1698 -299 -1690 -297
rect -1447 -311 -1439 -309
rect -1737 -323 -1729 -321
rect -1718 -323 -1710 -321
rect -1698 -323 -1690 -321
rect -1542 -326 -1534 -324
rect -1285 -326 -1277 -324
rect -1246 -326 -1238 -324
rect -1698 -351 -1690 -349
rect -1246 -350 -1238 -348
rect -2011 -359 -2003 -357
rect -1972 -359 -1964 -357
rect -1285 -362 -1277 -360
rect -1793 -366 -1785 -364
rect -1246 -374 -1238 -372
rect -1972 -383 -1964 -381
rect -2011 -395 -2003 -393
rect -1246 -398 -1238 -396
rect -1972 -407 -1964 -405
rect -1285 -422 -1277 -420
rect -1246 -422 -1238 -420
rect -1972 -431 -1964 -429
rect -1246 -446 -1238 -444
rect -2011 -455 -2003 -453
rect -1972 -455 -1964 -453
rect -1522 -456 -1514 -454
rect -1463 -457 -1455 -455
rect -1285 -470 -1277 -468
rect -1266 -470 -1258 -468
rect -1246 -470 -1238 -468
rect -1972 -479 -1964 -477
rect -1744 -479 -1736 -477
rect -1705 -479 -1697 -477
rect -2011 -503 -2003 -501
rect -1992 -503 -1984 -501
rect -1972 -503 -1964 -501
rect -1705 -503 -1697 -501
rect -1595 -483 -1587 -481
rect -1246 -498 -1238 -496
rect -1490 -500 -1482 -498
rect -1464 -500 -1456 -498
rect -1595 -505 -1587 -503
rect -1744 -515 -1736 -513
rect -1595 -524 -1587 -522
rect -1705 -527 -1697 -525
rect -1972 -531 -1964 -529
rect -2067 -546 -2059 -544
rect -1705 -551 -1697 -549
rect -1341 -513 -1333 -511
rect -1490 -534 -1482 -532
rect -1464 -534 -1456 -532
rect -1744 -575 -1736 -573
rect -1705 -575 -1697 -573
rect -1705 -599 -1697 -597
rect -1744 -623 -1736 -621
rect -1725 -623 -1717 -621
rect -1705 -623 -1697 -621
rect -1705 -651 -1697 -649
rect -1800 -666 -1792 -664
<< polycontact >>
rect -2056 222 -2052 226
rect -2031 221 -2027 225
rect -1967 221 -1963 225
rect -1942 220 -1938 224
rect -1880 221 -1876 225
rect -1855 220 -1851 224
rect -1791 222 -1787 226
rect -1766 221 -1762 225
rect -1703 222 -1699 226
rect -1678 221 -1674 225
rect -1613 222 -1609 226
rect -1588 221 -1584 225
rect -1521 222 -1517 226
rect -1496 221 -1492 225
rect -1426 222 -1422 226
rect -1401 221 -1397 225
rect -1337 222 -1333 226
rect -1312 221 -1308 225
rect -1245 223 -1241 227
rect -1220 222 -1216 226
rect -1151 222 -1147 226
rect -1126 221 -1122 225
rect -1063 222 -1059 226
rect -1038 221 -1034 225
rect -973 222 -969 226
rect -948 221 -944 225
rect -882 222 -878 226
rect -857 221 -853 225
rect -791 222 -787 226
rect -766 221 -762 225
rect -702 222 -698 226
rect -677 221 -673 225
rect -2028 180 -2024 184
rect -1939 179 -1935 183
rect -1852 179 -1848 183
rect -1763 180 -1759 184
rect -1675 180 -1671 184
rect -1585 180 -1581 184
rect -1493 180 -1489 184
rect -1398 180 -1394 184
rect -1309 180 -1305 184
rect -1217 181 -1213 185
rect -1123 180 -1119 184
rect -1035 180 -1031 184
rect -945 180 -941 184
rect -854 180 -850 184
rect -763 180 -759 184
rect -674 180 -670 184
rect -1955 73 -1951 77
rect -2000 63 -1996 67
rect -839 66 -835 70
rect -780 65 -776 69
rect -1962 39 -1958 43
rect -1703 43 -1699 47
rect -1644 42 -1640 46
rect -938 40 -934 44
rect -913 39 -909 43
rect -1287 33 -1283 37
rect -2014 27 -2010 31
rect -1228 32 -1224 36
rect -1992 15 -1988 19
rect -1802 17 -1798 21
rect -1777 16 -1773 20
rect -2243 -5 -2239 -1
rect -2288 -15 -2284 -11
rect -2044 -9 -2040 -5
rect -1705 10 -1701 14
rect -1386 7 -1382 11
rect -1361 6 -1357 10
rect -841 33 -837 37
rect -1774 -25 -1770 -21
rect -2016 -33 -2012 -29
rect -2006 -33 -2002 -29
rect -1951 -33 -1947 -29
rect -2250 -39 -2246 -35
rect -2302 -51 -2298 -47
rect -1969 -57 -1965 -53
rect -2280 -63 -2276 -59
rect -1644 -26 -1640 -22
rect -1289 0 -1285 4
rect -910 -2 -906 2
rect -1358 -35 -1354 -31
rect -1692 -47 -1688 -43
rect -1634 -64 -1630 -60
rect -1962 -71 -1958 -67
rect -2020 -81 -2016 -77
rect -1228 -36 -1224 -32
rect -780 -3 -776 1
rect -828 -24 -824 -20
rect -770 -41 -766 -37
rect -1276 -57 -1272 -53
rect -1218 -74 -1214 -70
rect -1043 -78 -1039 -74
rect -2332 -87 -2328 -83
rect -1088 -88 -1084 -84
rect -1962 -95 -1958 -91
rect -2304 -111 -2300 -107
rect -2294 -111 -2290 -107
rect -2239 -111 -2235 -107
rect -1957 -109 -1953 -105
rect -1050 -112 -1046 -108
rect -2052 -124 -2048 -120
rect -2257 -135 -2253 -131
rect -1461 -127 -1457 -123
rect -1102 -124 -1098 -120
rect -1506 -137 -1502 -133
rect -1080 -136 -1076 -132
rect -2250 -149 -2246 -145
rect -2308 -159 -2304 -155
rect -1468 -161 -1464 -157
rect -1132 -160 -1128 -156
rect -1712 -167 -1708 -163
rect -2250 -173 -2246 -169
rect -1757 -177 -1753 -173
rect -1520 -173 -1516 -169
rect -2245 -187 -2241 -183
rect -1498 -185 -1494 -181
rect -1104 -184 -1100 -180
rect -1094 -184 -1090 -180
rect -1039 -184 -1035 -180
rect -2340 -202 -2336 -198
rect -1719 -201 -1715 -197
rect -1771 -213 -1767 -209
rect -1550 -209 -1546 -205
rect -1057 -208 -1053 -204
rect -1749 -225 -1745 -221
rect -1050 -222 -1046 -218
rect -1522 -233 -1518 -229
rect -1512 -233 -1508 -229
rect -1457 -233 -1453 -229
rect -1108 -232 -1104 -228
rect -1801 -249 -1797 -245
rect -1050 -246 -1046 -242
rect -1475 -257 -1471 -253
rect -1045 -260 -1041 -256
rect -1773 -273 -1769 -269
rect -1763 -273 -1759 -269
rect -1708 -273 -1704 -269
rect -1468 -271 -1464 -267
rect -1526 -281 -1522 -277
rect -1140 -275 -1136 -271
rect -1726 -297 -1722 -293
rect -1468 -295 -1464 -291
rect -1719 -311 -1715 -307
rect -1463 -309 -1459 -305
rect -1777 -321 -1773 -317
rect -1260 -314 -1256 -310
rect -1558 -324 -1554 -320
rect -1305 -324 -1301 -320
rect -1719 -335 -1715 -331
rect -1986 -347 -1982 -343
rect -1714 -349 -1710 -345
rect -1267 -348 -1263 -344
rect -2031 -357 -2027 -353
rect -1809 -364 -1805 -360
rect -1319 -360 -1315 -356
rect -1297 -372 -1293 -368
rect -1993 -381 -1989 -377
rect -2045 -393 -2041 -389
rect -1349 -396 -1345 -392
rect -2023 -405 -2019 -401
rect -1321 -420 -1317 -416
rect -1311 -420 -1307 -416
rect -1256 -420 -1252 -416
rect -2075 -429 -2071 -425
rect -1274 -444 -1270 -440
rect -2047 -453 -2043 -449
rect -2037 -453 -2033 -449
rect -1982 -453 -1978 -449
rect -1535 -454 -1531 -450
rect -1476 -455 -1472 -451
rect -1267 -458 -1263 -454
rect -1719 -467 -1715 -463
rect -1325 -468 -1321 -464
rect -2000 -477 -1996 -473
rect -1764 -477 -1760 -473
rect -1634 -480 -1630 -476
rect -1609 -481 -1605 -477
rect -1993 -491 -1989 -487
rect -2051 -501 -2047 -497
rect -1726 -501 -1722 -497
rect -1993 -515 -1989 -511
rect -1778 -513 -1774 -509
rect -1267 -482 -1263 -478
rect -1537 -487 -1533 -483
rect -1262 -496 -1258 -492
rect -1988 -529 -1984 -525
rect -1756 -525 -1752 -521
rect -1606 -522 -1602 -518
rect -2083 -544 -2079 -540
rect -1808 -549 -1804 -545
rect -1476 -523 -1472 -519
rect -1357 -511 -1353 -507
rect -1524 -544 -1520 -540
rect -1466 -561 -1462 -557
rect -1780 -573 -1776 -569
rect -1770 -573 -1766 -569
rect -1715 -573 -1711 -569
rect -1733 -597 -1729 -593
rect -1726 -611 -1722 -607
rect -1784 -621 -1780 -617
rect -1726 -635 -1722 -631
rect -1721 -649 -1717 -645
rect -1816 -664 -1812 -660
<< ndcontact >>
rect -2060 210 -2056 214
rect -2043 210 -2039 214
rect -2060 202 -2056 206
rect -2043 202 -2039 206
rect -1971 209 -1967 213
rect -1954 209 -1950 213
rect -1971 201 -1967 205
rect -1954 201 -1950 205
rect -1884 209 -1880 213
rect -1867 209 -1863 213
rect -1884 201 -1880 205
rect -1867 201 -1863 205
rect -1795 210 -1791 214
rect -1778 210 -1774 214
rect -1795 202 -1791 206
rect -1778 202 -1774 206
rect -1707 210 -1703 214
rect -1690 210 -1686 214
rect -1707 202 -1703 206
rect -1690 202 -1686 206
rect -1617 210 -1613 214
rect -1600 210 -1596 214
rect -1617 202 -1613 206
rect -1600 202 -1596 206
rect -1525 210 -1521 214
rect -1508 210 -1504 214
rect -1525 202 -1521 206
rect -1508 202 -1504 206
rect -1430 210 -1426 214
rect -1413 210 -1409 214
rect -1430 202 -1426 206
rect -1413 202 -1409 206
rect -1341 210 -1337 214
rect -1324 210 -1320 214
rect -1341 202 -1337 206
rect -1324 202 -1320 206
rect -1249 211 -1245 215
rect -1232 211 -1228 215
rect -1249 203 -1245 207
rect -1232 203 -1228 207
rect -1155 210 -1151 214
rect -1138 210 -1134 214
rect -1155 202 -1151 206
rect -1138 202 -1134 206
rect -1067 210 -1063 214
rect -1050 210 -1046 214
rect -1067 202 -1063 206
rect -1050 202 -1046 206
rect -977 210 -973 214
rect -960 210 -956 214
rect -977 202 -973 206
rect -960 202 -956 206
rect -886 210 -882 214
rect -869 210 -865 214
rect -886 202 -882 206
rect -869 202 -865 206
rect -795 210 -791 214
rect -778 210 -774 214
rect -795 202 -791 206
rect -778 202 -774 206
rect -706 210 -702 214
rect -689 210 -685 214
rect -706 202 -702 206
rect -689 202 -685 206
rect -2042 181 -2038 185
rect -1953 180 -1949 184
rect -1866 180 -1862 184
rect -1777 181 -1773 185
rect -1689 181 -1685 185
rect -1599 181 -1595 185
rect -1507 181 -1503 185
rect -1412 181 -1408 185
rect -1323 181 -1319 185
rect -1231 182 -1227 186
rect -1137 181 -1133 185
rect -2042 173 -2038 177
rect -1049 181 -1045 185
rect -959 181 -955 185
rect -868 181 -864 185
rect -777 181 -773 185
rect -688 181 -684 185
rect -1953 172 -1949 176
rect -1866 172 -1862 176
rect -1777 173 -1773 177
rect -1689 173 -1685 177
rect -1599 173 -1595 177
rect -1507 173 -1503 177
rect -1412 173 -1408 177
rect -1323 173 -1319 177
rect -1231 174 -1227 178
rect -1137 173 -1133 177
rect -1049 173 -1045 177
rect -959 173 -955 177
rect -868 173 -864 177
rect -777 173 -773 177
rect -688 173 -684 177
rect -2061 64 -2057 68
rect -2028 64 -2024 68
rect -848 67 -844 71
rect -2061 56 -2057 60
rect -2028 56 -2024 60
rect -848 59 -844 63
rect -789 58 -785 62
rect -1712 44 -1708 48
rect -2061 40 -2057 44
rect -2061 32 -2057 36
rect -1712 36 -1708 40
rect -1653 35 -1649 39
rect -1296 34 -1292 38
rect -2028 28 -2024 32
rect -1296 26 -1292 30
rect -1237 25 -1233 29
rect -2028 20 -2024 24
rect -2061 16 -2057 20
rect -2061 8 -2057 12
rect -2349 -14 -2345 -10
rect -2316 -14 -2312 -10
rect -2061 -8 -2057 -4
rect -2061 -16 -2057 -12
rect -1806 5 -1802 9
rect -1789 5 -1785 9
rect -1806 -3 -1802 1
rect -1789 -3 -1785 1
rect -1709 -1 -1705 3
rect -1687 0 -1683 4
rect -942 28 -938 32
rect -925 28 -921 32
rect -942 20 -938 24
rect -925 20 -921 24
rect -845 22 -841 26
rect -823 23 -819 27
rect -845 14 -841 18
rect -1709 -9 -1705 -5
rect -2349 -22 -2345 -18
rect -2316 -22 -2312 -18
rect -1687 -8 -1683 -4
rect -1788 -24 -1784 -20
rect -2061 -32 -2057 -28
rect -2028 -32 -2024 -28
rect -1788 -32 -1784 -28
rect -2349 -38 -2345 -34
rect -2061 -40 -2057 -36
rect -2349 -46 -2345 -42
rect -2028 -40 -2024 -36
rect -2316 -50 -2312 -46
rect -2316 -58 -2312 -54
rect -2061 -56 -2057 -52
rect -2349 -62 -2345 -58
rect -2061 -64 -2057 -60
rect -2349 -70 -2345 -66
rect -1709 -28 -1705 -24
rect -1687 -27 -1683 -23
rect -1390 -5 -1386 -1
rect -823 15 -819 19
rect -1373 -5 -1369 -1
rect -1390 -13 -1386 -9
rect -1373 -13 -1369 -9
rect -1293 -11 -1289 -7
rect -1271 -10 -1267 -6
rect -924 -1 -920 3
rect -924 -9 -920 -5
rect -1293 -19 -1289 -15
rect -1271 -18 -1267 -14
rect -1709 -36 -1705 -32
rect -1687 -35 -1683 -31
rect -1372 -34 -1368 -30
rect -1372 -42 -1368 -38
rect -2061 -80 -2057 -76
rect -2044 -80 -2040 -76
rect -2028 -80 -2024 -76
rect -1293 -38 -1289 -34
rect -1271 -37 -1267 -33
rect -1293 -46 -1289 -42
rect -1271 -45 -1267 -41
rect -845 -5 -841 -1
rect -823 -4 -819 0
rect -845 -13 -841 -9
rect -823 -12 -819 -8
rect -2349 -86 -2345 -82
rect -2061 -88 -2057 -84
rect -2044 -88 -2040 -84
rect -2349 -94 -2345 -90
rect -2028 -88 -2024 -84
rect -1149 -87 -1145 -83
rect -1116 -87 -1112 -83
rect -1149 -95 -1145 -91
rect -1116 -95 -1112 -91
rect -2349 -110 -2345 -106
rect -2316 -110 -2312 -106
rect -1968 -108 -1964 -104
rect -1149 -111 -1145 -107
rect -2349 -118 -2345 -114
rect -2316 -118 -2312 -114
rect -1968 -116 -1964 -112
rect -1149 -119 -1145 -115
rect -2061 -123 -2057 -119
rect -1116 -123 -1112 -119
rect -2349 -134 -2345 -130
rect -2061 -131 -2057 -127
rect -1567 -136 -1563 -132
rect -1534 -136 -1530 -132
rect -1116 -131 -1112 -127
rect -1149 -135 -1145 -131
rect -2349 -142 -2345 -138
rect -1567 -144 -1563 -140
rect -1534 -144 -1530 -140
rect -1149 -143 -1145 -139
rect -2349 -158 -2345 -154
rect -2332 -158 -2328 -154
rect -2316 -158 -2312 -154
rect -1567 -160 -1563 -156
rect -1149 -159 -1145 -155
rect -2349 -166 -2345 -162
rect -2332 -166 -2328 -162
rect -2316 -166 -2312 -162
rect -1567 -168 -1563 -164
rect -1149 -167 -1145 -163
rect -1818 -176 -1814 -172
rect -1785 -176 -1781 -172
rect -1534 -172 -1530 -168
rect -2256 -186 -2252 -182
rect -1818 -184 -1814 -180
rect -1785 -184 -1781 -180
rect -1534 -180 -1530 -176
rect -1567 -184 -1563 -180
rect -1149 -183 -1145 -179
rect -1116 -183 -1112 -179
rect -2256 -194 -2252 -190
rect -1567 -192 -1563 -188
rect -1149 -191 -1145 -187
rect -1116 -191 -1112 -187
rect -2349 -201 -2345 -197
rect -1818 -200 -1814 -196
rect -2349 -209 -2345 -205
rect -1818 -208 -1814 -204
rect -1567 -208 -1563 -204
rect -1785 -212 -1781 -208
rect -1149 -207 -1145 -203
rect -1785 -220 -1781 -216
rect -1567 -216 -1563 -212
rect -1149 -215 -1145 -211
rect -1818 -224 -1814 -220
rect -1818 -232 -1814 -228
rect -1567 -232 -1563 -228
rect -1534 -232 -1530 -228
rect -1149 -231 -1145 -227
rect -1132 -231 -1128 -227
rect -1116 -231 -1112 -227
rect -1567 -240 -1563 -236
rect -1534 -240 -1530 -236
rect -1149 -239 -1145 -235
rect -1132 -239 -1128 -235
rect -1818 -248 -1814 -244
rect -1116 -239 -1112 -235
rect -1818 -256 -1814 -252
rect -1567 -256 -1563 -252
rect -1056 -259 -1052 -255
rect -1567 -264 -1563 -260
rect -1056 -267 -1052 -263
rect -1818 -272 -1814 -268
rect -1785 -272 -1781 -268
rect -1818 -280 -1814 -276
rect -1785 -280 -1781 -276
rect -1567 -280 -1563 -276
rect -1550 -280 -1546 -276
rect -1534 -280 -1530 -276
rect -1149 -274 -1145 -270
rect -1149 -282 -1145 -278
rect -1567 -288 -1563 -284
rect -1550 -288 -1546 -284
rect -1818 -296 -1814 -292
rect -1534 -288 -1530 -284
rect -1818 -304 -1814 -300
rect -1474 -308 -1470 -304
rect -1818 -320 -1814 -316
rect -1801 -320 -1797 -316
rect -1785 -320 -1781 -316
rect -1474 -316 -1470 -312
rect -1567 -323 -1563 -319
rect -1818 -328 -1814 -324
rect -1801 -328 -1797 -324
rect -1785 -328 -1781 -324
rect -1366 -323 -1362 -319
rect -1333 -323 -1329 -319
rect -1567 -331 -1563 -327
rect -1366 -331 -1362 -327
rect -1333 -331 -1329 -327
rect -1725 -348 -1721 -344
rect -1366 -347 -1362 -343
rect -2092 -356 -2088 -352
rect -2059 -356 -2055 -352
rect -1725 -356 -1721 -352
rect -1366 -355 -1362 -351
rect -1333 -359 -1329 -355
rect -2092 -364 -2088 -360
rect -2059 -364 -2055 -360
rect -1818 -363 -1814 -359
rect -1818 -371 -1814 -367
rect -1333 -367 -1329 -363
rect -1366 -371 -1362 -367
rect -2092 -380 -2088 -376
rect -1366 -379 -1362 -375
rect -2092 -388 -2088 -384
rect -2059 -392 -2055 -388
rect -1366 -395 -1362 -391
rect -2059 -400 -2055 -396
rect -2092 -404 -2088 -400
rect -1366 -403 -1362 -399
rect -2092 -412 -2088 -408
rect -1366 -419 -1362 -415
rect -1333 -419 -1329 -415
rect -2092 -428 -2088 -424
rect -1366 -427 -1362 -423
rect -1333 -427 -1329 -423
rect -2092 -436 -2088 -432
rect -1366 -443 -1362 -439
rect -2092 -452 -2088 -448
rect -2059 -452 -2055 -448
rect -1544 -453 -1540 -449
rect -2092 -460 -2088 -456
rect -2059 -460 -2055 -456
rect -1366 -451 -1362 -447
rect -1544 -461 -1540 -457
rect -1485 -462 -1481 -458
rect -1366 -467 -1362 -463
rect -1349 -467 -1345 -463
rect -1333 -467 -1329 -463
rect -2092 -476 -2088 -472
rect -1825 -476 -1821 -472
rect -1792 -476 -1788 -472
rect -1366 -475 -1362 -471
rect -1349 -475 -1345 -471
rect -2092 -484 -2088 -480
rect -1825 -484 -1821 -480
rect -1792 -484 -1788 -480
rect -1333 -475 -1329 -471
rect -2092 -500 -2088 -496
rect -2075 -500 -2071 -496
rect -2059 -500 -2055 -496
rect -1825 -500 -1821 -496
rect -2092 -508 -2088 -504
rect -2075 -508 -2071 -504
rect -2059 -508 -2055 -504
rect -1825 -508 -1821 -504
rect -1792 -512 -1788 -508
rect -1638 -492 -1634 -488
rect -1621 -492 -1617 -488
rect -1638 -500 -1634 -496
rect -1621 -500 -1617 -496
rect -1541 -498 -1537 -494
rect -1519 -497 -1515 -493
rect -1273 -495 -1269 -491
rect -1541 -506 -1537 -502
rect -1519 -505 -1515 -501
rect -1792 -520 -1788 -516
rect -1825 -524 -1821 -520
rect -1999 -528 -1995 -524
rect -1620 -521 -1616 -517
rect -1999 -536 -1995 -532
rect -1825 -532 -1821 -528
rect -1620 -529 -1616 -525
rect -2092 -543 -2088 -539
rect -2092 -551 -2088 -547
rect -1825 -548 -1821 -544
rect -1825 -556 -1821 -552
rect -1541 -525 -1537 -521
rect -1519 -524 -1515 -520
rect -1273 -503 -1269 -499
rect -1366 -510 -1362 -506
rect -1366 -518 -1362 -514
rect -1541 -533 -1537 -529
rect -1519 -532 -1515 -528
rect -1825 -572 -1821 -568
rect -1792 -572 -1788 -568
rect -1825 -580 -1821 -576
rect -1792 -580 -1788 -576
rect -1825 -596 -1821 -592
rect -1825 -604 -1821 -600
rect -1825 -620 -1821 -616
rect -1808 -620 -1804 -616
rect -1792 -620 -1788 -616
rect -1825 -628 -1821 -624
rect -1808 -628 -1804 -624
rect -1792 -628 -1788 -624
rect -1732 -648 -1728 -644
rect -1732 -656 -1728 -652
rect -1825 -663 -1821 -659
rect -1825 -671 -1821 -667
<< pdcontact >>
rect -2017 222 -2009 226
rect -1928 221 -1920 225
rect -2017 214 -2009 218
rect -2017 200 -2009 204
rect -2017 192 -2009 196
rect -1841 221 -1833 225
rect -1752 222 -1744 226
rect -1928 213 -1920 217
rect -1928 199 -1920 203
rect -1928 191 -1920 195
rect -1841 213 -1833 217
rect -1841 199 -1833 203
rect -1841 191 -1833 195
rect -1664 222 -1656 226
rect -1752 214 -1744 218
rect -1752 200 -1744 204
rect -1752 192 -1744 196
rect -1574 222 -1566 226
rect -1664 214 -1656 218
rect -1664 200 -1656 204
rect -1664 192 -1656 196
rect -1482 222 -1474 226
rect -1574 214 -1566 218
rect -1574 200 -1566 204
rect -1574 192 -1566 196
rect -1387 222 -1379 226
rect -1482 214 -1474 218
rect -1482 200 -1474 204
rect -1482 192 -1474 196
rect -1298 222 -1290 226
rect -1206 223 -1198 227
rect -1387 214 -1379 218
rect -1387 200 -1379 204
rect -1387 192 -1379 196
rect -1298 214 -1290 218
rect -1298 200 -1290 204
rect -1298 192 -1290 196
rect -1112 222 -1104 226
rect -1206 215 -1198 219
rect -1206 201 -1198 205
rect -1206 193 -1198 197
rect -1024 222 -1016 226
rect -1112 214 -1104 218
rect -1112 200 -1104 204
rect -1112 192 -1104 196
rect -934 222 -926 226
rect -1024 214 -1016 218
rect -1024 200 -1016 204
rect -1024 192 -1016 196
rect -843 222 -835 226
rect -934 214 -926 218
rect -934 200 -926 204
rect -934 192 -926 196
rect -752 222 -744 226
rect -843 214 -835 218
rect -843 200 -835 204
rect -843 192 -835 196
rect -663 222 -655 226
rect -752 214 -744 218
rect -752 200 -744 204
rect -752 192 -744 196
rect -663 214 -655 218
rect -663 200 -655 204
rect -663 192 -655 196
rect -2017 181 -2009 185
rect -1928 180 -1920 184
rect -1841 180 -1833 184
rect -1752 181 -1744 185
rect -1664 181 -1656 185
rect -1574 181 -1566 185
rect -1482 181 -1474 185
rect -1387 181 -1379 185
rect -1298 181 -1290 185
rect -1206 182 -1198 186
rect -1112 181 -1104 185
rect -1024 181 -1016 185
rect -934 181 -926 185
rect -843 181 -835 185
rect -752 181 -744 185
rect -663 181 -655 185
rect -2017 173 -2009 177
rect -1928 172 -1920 176
rect -1841 172 -1833 176
rect -1752 173 -1744 177
rect -1664 173 -1656 177
rect -1574 173 -1566 177
rect -1482 173 -1474 177
rect -1387 173 -1379 177
rect -1298 173 -1290 177
rect -1206 174 -1199 178
rect -1112 173 -1104 177
rect -1024 173 -1016 177
rect -934 173 -926 177
rect -843 173 -835 177
rect -752 173 -744 177
rect -663 173 -655 177
rect -1980 64 -1972 68
rect -1941 64 -1933 68
rect -826 67 -818 71
rect -767 66 -759 70
rect -1980 56 -1972 60
rect -1941 56 -1933 60
rect -826 59 -818 63
rect -767 58 -759 62
rect -1941 40 -1933 44
rect -1690 44 -1682 48
rect -1631 43 -1623 47
rect -1690 36 -1682 40
rect -1941 32 -1933 36
rect -1631 35 -1623 39
rect -899 40 -891 44
rect -1274 34 -1266 38
rect -1980 28 -1972 32
rect -1215 33 -1207 37
rect -1274 26 -1266 30
rect -1215 25 -1207 29
rect -1980 20 -1972 24
rect -1941 16 -1933 20
rect -1763 17 -1755 21
rect -1941 8 -1933 12
rect -2268 -14 -2260 -10
rect -1941 -8 -1933 -4
rect -2229 -14 -2221 -10
rect -1941 -16 -1933 -12
rect -1763 9 -1755 13
rect -1763 -5 -1755 -1
rect -1347 7 -1339 11
rect -899 32 -891 36
rect -899 18 -891 22
rect -794 23 -786 27
rect -768 23 -760 27
rect -899 10 -891 14
rect -1658 0 -1650 4
rect -1632 0 -1624 4
rect -1763 -13 -1755 -9
rect -2268 -22 -2260 -18
rect -1658 -8 -1650 -4
rect -2229 -22 -2221 -18
rect -1763 -24 -1755 -20
rect -1980 -32 -1972 -28
rect -1941 -32 -1933 -28
rect -1763 -32 -1755 -28
rect -2229 -38 -2221 -34
rect -2229 -46 -2221 -42
rect -1980 -40 -1972 -36
rect -1941 -40 -1933 -36
rect -2268 -50 -2260 -46
rect -2268 -58 -2260 -54
rect -1941 -56 -1933 -52
rect -2229 -62 -2221 -58
rect -1941 -64 -1933 -60
rect -2229 -70 -2221 -66
rect -1632 -8 -1624 -4
rect -794 15 -786 19
rect -1347 -1 -1339 3
rect -1347 -15 -1339 -11
rect -899 -1 -891 3
rect -1242 -10 -1234 -6
rect -1216 -10 -1208 -6
rect -899 -9 -891 -5
rect -1347 -23 -1339 -19
rect -1242 -18 -1234 -14
rect -1658 -34 -1650 -30
rect -1632 -34 -1624 -30
rect -1347 -34 -1339 -30
rect -1658 -42 -1650 -38
rect -1632 -42 -1624 -38
rect -1347 -42 -1339 -38
rect -1980 -80 -1972 -76
rect -1961 -80 -1953 -76
rect -1216 -18 -1208 -14
rect -1242 -44 -1234 -40
rect -1216 -44 -1208 -40
rect -768 15 -760 19
rect -794 -11 -786 -7
rect -768 -11 -760 -7
rect -794 -19 -786 -15
rect -768 -19 -760 -15
rect -1242 -52 -1234 -48
rect -1216 -52 -1208 -48
rect -1941 -80 -1933 -76
rect -2229 -86 -2221 -82
rect -2229 -94 -2221 -90
rect -1980 -88 -1972 -84
rect -1961 -88 -1953 -84
rect -1941 -88 -1933 -84
rect -1068 -87 -1060 -83
rect -1029 -87 -1021 -83
rect -1068 -95 -1060 -91
rect -1029 -95 -1021 -91
rect -2268 -110 -2260 -106
rect -2229 -110 -2221 -106
rect -1941 -108 -1933 -104
rect -2268 -118 -2260 -114
rect -2229 -118 -2221 -114
rect -1029 -111 -1021 -107
rect -1941 -116 -1933 -112
rect -1029 -119 -1021 -115
rect -2036 -123 -2028 -119
rect -2229 -134 -2221 -130
rect -1068 -123 -1060 -119
rect -2036 -131 -2028 -127
rect -1486 -136 -1478 -132
rect -1068 -131 -1060 -127
rect -1447 -136 -1439 -132
rect -1029 -135 -1021 -131
rect -2229 -142 -2221 -138
rect -1486 -144 -1478 -140
rect -1447 -144 -1439 -140
rect -1029 -143 -1021 -139
rect -2268 -158 -2260 -154
rect -2249 -158 -2241 -154
rect -2229 -158 -2221 -154
rect -1447 -160 -1439 -156
rect -1029 -159 -1021 -155
rect -2268 -166 -2260 -162
rect -2249 -166 -2241 -162
rect -2229 -166 -2221 -162
rect -1447 -168 -1439 -164
rect -1029 -167 -1021 -163
rect -1737 -176 -1729 -172
rect -1698 -176 -1690 -172
rect -1486 -172 -1478 -168
rect -2229 -186 -2221 -182
rect -1737 -184 -1729 -180
rect -1486 -180 -1478 -176
rect -1698 -184 -1690 -180
rect -1447 -184 -1439 -180
rect -1068 -183 -1060 -179
rect -1029 -183 -1021 -179
rect -2229 -194 -2221 -190
rect -1447 -192 -1439 -188
rect -1068 -191 -1060 -187
rect -1029 -191 -1021 -187
rect -2324 -201 -2316 -197
rect -1698 -200 -1690 -196
rect -2324 -209 -2316 -205
rect -1698 -208 -1690 -204
rect -1737 -212 -1729 -208
rect -1447 -208 -1439 -204
rect -1029 -207 -1021 -203
rect -1447 -216 -1439 -212
rect -1029 -215 -1021 -211
rect -1737 -220 -1729 -216
rect -1698 -224 -1690 -220
rect -1698 -232 -1690 -228
rect -1486 -232 -1478 -228
rect -1447 -232 -1439 -228
rect -1068 -231 -1060 -227
rect -1049 -231 -1041 -227
rect -1029 -231 -1021 -227
rect -1486 -240 -1478 -236
rect -1447 -240 -1439 -236
rect -1698 -248 -1690 -244
rect -1068 -239 -1060 -235
rect -1049 -239 -1041 -235
rect -1029 -239 -1021 -235
rect -1698 -256 -1690 -252
rect -1447 -256 -1439 -252
rect -1029 -259 -1021 -255
rect -1447 -264 -1439 -260
rect -1029 -267 -1021 -263
rect -1737 -272 -1729 -268
rect -1698 -272 -1690 -268
rect -1737 -280 -1729 -276
rect -1698 -280 -1690 -276
rect -1486 -280 -1478 -276
rect -1467 -280 -1459 -276
rect -1124 -274 -1116 -270
rect -1447 -280 -1439 -276
rect -1124 -282 -1116 -278
rect -1698 -296 -1690 -292
rect -1486 -288 -1478 -284
rect -1467 -288 -1459 -284
rect -1447 -288 -1439 -284
rect -1698 -304 -1690 -300
rect -1447 -308 -1439 -304
rect -1737 -320 -1729 -316
rect -1718 -320 -1710 -316
rect -1447 -316 -1439 -312
rect -1698 -320 -1690 -316
rect -1737 -328 -1729 -324
rect -1718 -328 -1710 -324
rect -1542 -323 -1534 -319
rect -1285 -323 -1277 -319
rect -1246 -323 -1238 -319
rect -1698 -328 -1690 -324
rect -1542 -331 -1534 -327
rect -1285 -331 -1277 -327
rect -1246 -331 -1238 -327
rect -1698 -348 -1690 -344
rect -1246 -347 -1238 -343
rect -2011 -356 -2003 -352
rect -1972 -356 -1964 -352
rect -1698 -356 -1690 -352
rect -1246 -355 -1238 -351
rect -2011 -364 -2003 -360
rect -1972 -364 -1964 -360
rect -1793 -363 -1785 -359
rect -1285 -359 -1277 -355
rect -1285 -367 -1277 -363
rect -1793 -371 -1785 -367
rect -1246 -371 -1238 -367
rect -1972 -380 -1964 -376
rect -1246 -379 -1238 -375
rect -1972 -388 -1964 -384
rect -2011 -392 -2003 -388
rect -1246 -395 -1238 -391
rect -2011 -400 -2003 -396
rect -1972 -404 -1964 -400
rect -1246 -403 -1238 -399
rect -1972 -412 -1964 -408
rect -1285 -419 -1277 -415
rect -1246 -419 -1238 -415
rect -1972 -428 -1964 -424
rect -1285 -427 -1277 -423
rect -1246 -427 -1238 -423
rect -1972 -436 -1964 -432
rect -1246 -443 -1238 -439
rect -2011 -452 -2003 -448
rect -1972 -452 -1964 -448
rect -1522 -453 -1514 -449
rect -2011 -460 -2003 -456
rect -1463 -454 -1455 -450
rect -1246 -451 -1238 -447
rect -1972 -460 -1964 -456
rect -1522 -461 -1514 -457
rect -1463 -462 -1455 -458
rect -1285 -467 -1277 -463
rect -1266 -467 -1258 -463
rect -1246 -467 -1238 -463
rect -1972 -476 -1964 -472
rect -1744 -476 -1736 -472
rect -1705 -476 -1697 -472
rect -1972 -484 -1964 -480
rect -1744 -484 -1736 -480
rect -1705 -484 -1697 -480
rect -1595 -480 -1587 -476
rect -1285 -475 -1277 -471
rect -1266 -475 -1258 -471
rect -1246 -475 -1238 -471
rect -2011 -500 -2003 -496
rect -1992 -500 -1984 -496
rect -1972 -500 -1964 -496
rect -1705 -500 -1697 -496
rect -2011 -508 -2003 -504
rect -1992 -508 -1984 -504
rect -1972 -508 -1964 -504
rect -1705 -508 -1697 -504
rect -1744 -512 -1736 -508
rect -1595 -488 -1587 -484
rect -1595 -502 -1587 -498
rect -1490 -497 -1482 -493
rect -1464 -497 -1456 -493
rect -1246 -495 -1238 -491
rect -1595 -510 -1587 -506
rect -1490 -505 -1482 -501
rect -1744 -520 -1736 -516
rect -1972 -528 -1964 -524
rect -1705 -524 -1697 -520
rect -1595 -521 -1587 -517
rect -1705 -532 -1697 -528
rect -1595 -529 -1587 -525
rect -1972 -536 -1964 -532
rect -2067 -543 -2059 -539
rect -2067 -551 -2059 -547
rect -1705 -548 -1697 -544
rect -1705 -556 -1697 -552
rect -1464 -505 -1456 -501
rect -1246 -503 -1238 -499
rect -1341 -510 -1333 -506
rect -1341 -518 -1333 -514
rect -1490 -531 -1482 -527
rect -1464 -531 -1456 -527
rect -1490 -539 -1482 -535
rect -1464 -539 -1456 -535
rect -1744 -572 -1736 -568
rect -1705 -572 -1697 -568
rect -1744 -580 -1736 -576
rect -1705 -580 -1697 -576
rect -1705 -596 -1697 -592
rect -1705 -604 -1697 -600
rect -1744 -620 -1736 -616
rect -1725 -620 -1717 -616
rect -1705 -620 -1697 -616
rect -1744 -628 -1736 -624
rect -1725 -628 -1717 -624
rect -1705 -628 -1697 -624
rect -1705 -648 -1697 -644
rect -1705 -656 -1697 -652
rect -1800 -663 -1792 -659
rect -1800 -671 -1792 -667
<< m2contact >>
rect -1814 242 -1810 246
rect -2332 -79 -2328 -75
rect -1828 133 -1824 137
rect -1838 109 -1834 113
rect -2044 -1 -2040 3
rect -2075 -421 -2071 -417
rect -1362 242 -1358 246
rect -1765 148 -1761 152
rect -1677 133 -1673 137
rect -907 242 -903 246
rect -1362 150 -1358 154
rect -1781 109 -1777 113
rect -1802 94 -1798 98
rect -1419 127 -1414 131
rect -1644 94 -1640 98
rect -1814 5 -1810 9
rect -1747 -39 -1741 -33
rect -1747 -83 -1741 -78
rect -1141 100 -1137 104
rect -1386 84 -1382 88
rect -1398 80 -1394 84
rect -1066 100 -1062 104
rect -1228 84 -1224 88
rect -1398 -5 -1394 -1
rect -1419 -81 -1414 -77
rect -1419 -98 -1414 -94
rect -1331 -49 -1325 -43
rect -1331 -93 -1325 -88
rect -1801 -241 -1797 -237
rect -1419 -118 -1414 -114
rect -938 117 -934 121
rect -780 117 -776 121
rect -950 28 -946 32
rect -883 -16 -877 -10
rect -883 -60 -877 -55
rect -1550 -201 -1546 -197
rect -1578 -323 -1574 -319
rect -1848 -417 -1844 -413
rect -1664 -450 -1660 -446
rect -1132 -152 -1128 -148
rect -1557 -355 -1552 -351
rect -1349 -388 -1345 -384
rect -1535 -394 -1531 -390
rect -1634 -403 -1630 -399
rect -1476 -403 -1472 -399
rect -1646 -492 -1642 -488
rect -1808 -541 -1804 -537
rect -1579 -536 -1573 -530
rect -1579 -580 -1573 -575
rect -1721 -688 -1717 -684
<< labels >>
rlabel metal1 -677 246 -673 250 5 A0
rlabel metal1 -702 246 -698 250 5 B0
rlabel metal1 -676 -570 -672 -566 1 P0
rlabel metal2 -647 159 -641 163 7 n1
rlabel metal2 -714 242 -710 246 1 gnd
rlabel space -959 -103 -720 150 3 HalfAdder
rlabel metal1 -2339 -234 -2334 -230 1 CO
rlabel metal1 -2245 -226 -2241 -222 1 P6
rlabel metal1 -1510 -640 -1505 -636 1 P4
rlabel metal1 -1262 -635 -1258 -631 1 P3
rlabel metal1 -1045 -560 -1041 -556 1 P2
rlabel metal1 -814 -570 -809 -566 1 P1
rlabel metal1 -2056 246 -2052 250 5 B3
rlabel metal1 -2031 246 -2027 250 5 A3
rlabel space -1967 246 -1963 250 5 B2
rlabel space -1942 246 -1938 250 5 A3
rlabel space -1880 246 -1876 250 5 A2
rlabel space -1855 246 -1851 250 5 B3
rlabel metal1 -1791 246 -1787 250 5 B3
rlabel metal1 -1766 246 -1762 250 5 A1
rlabel metal1 -1703 246 -1699 250 5 A3
rlabel metal1 -1678 246 -1674 250 5 B1
rlabel metal1 -1613 246 -1609 250 5 B2
rlabel metal1 -1588 246 -1584 250 5 A2
rlabel metal1 -1521 246 -1517 250 5 A2
rlabel metal1 -1496 246 -1492 250 5 B1
rlabel metal1 -1426 246 -1422 250 5 B0
rlabel metal1 -1401 246 -1397 250 5 A3
rlabel metal1 -1337 246 -1333 250 5 A0
rlabel metal1 -1312 246 -1308 250 5 B3
rlabel metal1 -1245 247 -1241 251 5 B2
rlabel metal1 -1220 247 -1216 251 5 A1
rlabel metal1 -1151 246 -1147 250 5 B1
rlabel space -1126 247 -1122 251 5 A1
rlabel metal1 -1063 246 -1059 250 5 A2
rlabel metal1 -1038 246 -1034 250 5 B0
rlabel metal1 -973 246 -969 250 5 B2
rlabel metal1 -948 246 -944 250 5 A0
rlabel metal1 -882 246 -878 250 5 A1
rlabel metal1 -857 246 -853 250 5 B0
rlabel metal1 -791 246 -787 250 5 B1
rlabel metal1 -766 246 -762 250 5 A0
rlabel space -1564 -580 -1430 -413 3 XOR
rlabel space -1732 -83 -1598 84 3 XOR
rlabel space -1316 -93 -1182 74 3 XOR
rlabel space -868 -60 -734 107 3 XOR
rlabel space -1427 -155 -1128 34 1 fulladder
rlabel metal1 -1988 -729 -1984 -725 1 P5
<< end >>
