module multiplier(a0,a1,a2,a3,b0,b1,b2,b3,p0,p1,p2,p3,p4,p5,p6,c);

    input a0;
    input a1;
    input a2;
    input a3;
    input b0;
    input b1;
    input b2;
    input b3;
    output p0;
    output p1;
    output p2;
    output p3;
    output p4;
    output p5;
    output p6;
    output c;

    and(p0,a0,b0);
    and(o0,a0,b1);
    and(o1,a1,b0);
    and(o2,b2,a0);
    and(o3,a2,b0);
    and(o4,a1,b1);
    and(o5,a1,b2);
    and(o6,a0,b3);
    and(o7,a3,b0);
    and(o8,a2,b1);
    and(o9,a2,b2);
    and(o10,a3,b1);
    and(o11,a1,b3);
    and(o12,a2,b3);
    and(o13,a3,b2);
    and(o14,a3,b3);

    xor(p1,o0,o1);
    and(c0,o0,o1);
    xor(s0,o3,o4);
    and(c2,o3,o4);
    xor(s1,o7,o8);
    and(c3,o7,o8);
    xor(p4,s4,c5);
    and(c8,s4,c5);

    xor(p2,c0,o2,s0);
    xor(y1,c0,o2);
    and(y2,c0,o2);
    and(y3,y1,s0);
    or(c1,y2,y3);
    xor(s2,s1,o5,c2);
    xor(y4,s1,o5);
    and(y5,s1,o5);
    and(y6,y4,s2);
    or(c4,y5,y6);
    xor(p3,o6,c1,s2);
    xor(y7,o6,c1);
    and(y8,o6,c1);
    and(y9,y7,s2);
    or(c5,y8,y9);
    xor(s3,c3,o9,o10);
    xor(y10,c3,o9);
    and(y11,c3,o9);
    and(y12,y10,o10);
    or(c6,y11,y12);
    xor(s4,s3,c4,o11);
    xor(y13,s3,c4);
    and(y14,s3,c4);
    and(y15,y13,o11);
    or(c7,y14,y15);
    xor(s5,o13,o12,c6);
    xor(y16,o13,o12);
    and(y17,o13,o12);
    and(y18,y16,c6);
    or(c9,y17,y18);
    xor(p5,c7,c8,s5);
    xor(y19,c7,c8);
    and(y20,c7,c8);
    and(y21,y19,s5);
    or(c10,y20,y21);
    xor(p6,o14,c9,c10);
    xor(y22,o14,c9);
    and(y23,o14,c9);
    and(y24,y22,c10);
    or(c,y23,y24);

endmodule